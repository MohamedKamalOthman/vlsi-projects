/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 16:04:24 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2881660147 */

module n_case(A, B, S, outA, outB, enable);
   input [31:0]A;
   input [31:0]B;
   output [31:0]S;
   output [2:0]outA;
   output [2:0]outB;
   output enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_4;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;

   AND2_X1 i_0_0 (.A1(outB[0]), .A2(outA[0]), .ZN(enable));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(S[22]));
   OAI22_X1 i_0_2 (.A1(outB[1]), .A2(outB[0]), .B1(outA[1]), .B2(outA[0]), 
      .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(S[30]));
   OAI22_X1 i_0_4 (.A1(n_0_21), .A2(outA[2]), .B1(n_0_16), .B2(outB[2]), 
      .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(S[31]));
   XNOR2_X1 i_0_6 (.A(B[31]), .B(A[31]), .ZN(n_0_2));
   AOI22_X1 i_0_7 (.A1(outA[2]), .A2(n_0_5), .B1(n_0_7), .B2(outB[2]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_21), .A2(n_0_17), .ZN(n_0_5));
   AOI21_X1 i_0_9 (.A(outA[2]), .B1(n_0_28), .B2(n_0_17), .ZN(outA[0]));
   AOI21_X1 i_0_10 (.A(n_0_28), .B1(n_0_17), .B2(outA[2]), .ZN(outA[1]));
   NOR2_X1 i_0_11 (.A1(n_0_20), .A2(n_0_19), .ZN(outA[2]));
   NAND4_X1 i_0_12 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_0_19));
   NAND4_X1 i_0_13 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(outB[2]), .B1(n_0_31), .B2(n_0_8), .ZN(outB[0]));
   NAND2_X1 i_0_15 (.A1(n_0_31), .A2(n_0_8), .ZN(n_0_21));
   AOI21_X1 i_0_16 (.A(n_0_31), .B1(n_0_8), .B2(outB[2]), .ZN(outB[1]));
   AND2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_32), .ZN(n_0_31));
   NOR4_X1 i_0_18 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_32));
   NOR4_X1 i_0_19 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_33));
   NOR2_X1 i_0_20 (.A1(n_0_6), .A2(n_0_4), .ZN(outB[2]));
   NAND4_X1 i_0_21 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_4));
   NAND4_X1 i_0_22 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_6));
   NAND2_X1 i_0_23 (.A1(n_0_16), .A2(n_0_8), .ZN(n_0_7));
   AND3_X1 i_0_24 (.A1(n_0_10), .A2(n_0_9), .A3(n_0_11), .ZN(n_0_8));
   NOR4_X1 i_0_25 (.A1(B[19]), .A2(B[18]), .A3(B[16]), .A4(B[12]), .ZN(n_0_9));
   NOR4_X1 i_0_26 (.A1(B[17]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n_0_10));
   NOR4_X1 i_0_27 (.A1(B[10]), .A2(B[9]), .A3(B[8]), .A4(n_0_12), .ZN(n_0_11));
   NAND3_X1 i_0_28 (.A1(n_0_14), .A2(n_0_13), .A3(n_0_15), .ZN(n_0_12));
   NOR4_X1 i_0_29 (.A1(B[5]), .A2(B[3]), .A3(B[2]), .A4(B[1]), .ZN(n_0_13));
   NOR4_X1 i_0_30 (.A1(B[22]), .A2(B[21]), .A3(B[20]), .A4(B[0]), .ZN(n_0_14));
   NOR4_X1 i_0_31 (.A1(B[11]), .A2(B[7]), .A3(B[6]), .A4(B[4]), .ZN(n_0_15));
   NAND2_X1 i_0_32 (.A1(n_0_28), .A2(n_0_17), .ZN(n_0_16));
   AND3_X1 i_0_33 (.A1(n_0_22), .A2(n_0_18), .A3(n_0_23), .ZN(n_0_17));
   NOR4_X1 i_0_34 (.A1(A[19]), .A2(A[18]), .A3(A[16]), .A4(A[12]), .ZN(n_0_18));
   NOR4_X1 i_0_35 (.A1(A[17]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n_0_22));
   NOR4_X1 i_0_36 (.A1(A[10]), .A2(A[9]), .A3(A[8]), .A4(n_0_24), .ZN(n_0_23));
   NAND3_X1 i_0_37 (.A1(n_0_26), .A2(n_0_25), .A3(n_0_27), .ZN(n_0_24));
   NOR4_X1 i_0_38 (.A1(A[5]), .A2(A[3]), .A3(A[2]), .A4(A[1]), .ZN(n_0_25));
   NOR4_X1 i_0_39 (.A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[0]), .ZN(n_0_26));
   NOR4_X1 i_0_40 (.A1(A[11]), .A2(A[7]), .A3(A[6]), .A4(A[4]), .ZN(n_0_27));
   AND2_X1 i_0_41 (.A1(n_0_30), .A2(n_0_29), .ZN(n_0_28));
   NOR4_X1 i_0_42 (.A1(A[25]), .A2(A[24]), .A3(A[30]), .A4(A[27]), .ZN(n_0_29));
   NOR4_X1 i_0_43 (.A1(A[26]), .A2(A[23]), .A3(A[29]), .A4(A[28]), .ZN(n_0_30));
endmodule

module zero_counter(M, Zcount);
   input [23:0]M;
   output [4:0]Zcount;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_0), .B2(Zcount[4]), .ZN(Zcount[0]));
   OAI21_X1 i_0_1 (.A(n_0_33), .B1(M[6]), .B2(n_0_1), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(M[5]), .A2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(M[4]), .A2(n_0_3), .ZN(n_0_2));
   NOR2_X1 i_0_4 (.A1(M[3]), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(M[2]), .B1(n_0_32), .B2(M[0]), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(n_0_6), .B1(n_0_9), .B2(n_0_27), .ZN(n_0_5));
   AOI211_X1 i_0_7 (.A(M[15]), .B(n_0_27), .C1(n_0_7), .C2(n_0_36), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_35), .B1(M[12]), .B2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(M[11]), .B1(n_0_34), .B2(M[9]), .ZN(n_0_8));
   AOI221_X1 i_0_10 (.A(M[23]), .B1(n_0_39), .B2(M[21]), .C1(n_0_30), .C2(n_0_10), 
      .ZN(n_0_9));
   OAI21_X1 i_0_11 (.A(n_0_38), .B1(n_0_37), .B2(M[18]), .ZN(n_0_10));
   AOI21_X1 i_0_12 (.A(n_0_14), .B1(n_0_11), .B2(Zcount[4]), .ZN(Zcount[1]));
   OR3_X1 i_0_13 (.A1(M[7]), .A2(M[6]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(M[5]), .A2(M[4]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(M[3]), .A2(M[2]), .A3(n_0_23), .ZN(n_0_13));
   AOI22_X1 i_0_16 (.A1(n_0_26), .A2(n_0_17), .B1(n_0_15), .B2(n_0_27), .ZN(
      n_0_14));
   NOR3_X1 i_0_17 (.A1(M[23]), .A2(M[22]), .A3(n_0_16), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(M[21]), .A2(M[20]), .A3(n_0_29), .ZN(n_0_16));
   OAI21_X1 i_0_19 (.A(n_0_25), .B1(M[10]), .B2(M[11]), .ZN(n_0_17));
   OAI21_X1 i_0_20 (.A(n_0_18), .B1(n_0_19), .B2(Zcount[4]), .ZN(Zcount[2]));
   NAND3_X1 i_0_21 (.A1(Zcount[4]), .A2(n_0_22), .A3(n_0_21), .ZN(n_0_18));
   AOI22_X1 i_0_22 (.A1(n_0_26), .A2(n_0_25), .B1(n_0_30), .B2(n_0_27), .ZN(
      n_0_19));
   OAI22_X1 i_0_23 (.A1(n_0_22), .A2(n_0_20), .B1(n_0_27), .B2(Zcount[4]), 
      .ZN(Zcount[3]));
   NAND2_X1 i_0_24 (.A1(Zcount[4]), .A2(n_0_21), .ZN(n_0_20));
   NOR4_X1 i_0_25 (.A1(M[7]), .A2(M[6]), .A3(M[5]), .A4(M[4]), .ZN(n_0_21));
   NAND2_X1 i_0_26 (.A1(n_0_24), .A2(n_0_23), .ZN(n_0_22));
   NOR2_X1 i_0_27 (.A1(M[1]), .A2(M[0]), .ZN(n_0_23));
   NOR2_X1 i_0_28 (.A1(M[3]), .A2(M[2]), .ZN(n_0_24));
   AND3_X1 i_0_29 (.A1(n_0_31), .A2(n_0_26), .A3(n_0_25), .ZN(Zcount[4]));
   NOR2_X1 i_0_30 (.A1(M[13]), .A2(M[12]), .ZN(n_0_25));
   NOR3_X1 i_0_31 (.A1(n_0_27), .A2(M[14]), .A3(M[15]), .ZN(n_0_26));
   NAND3_X1 i_0_32 (.A1(n_0_30), .A2(n_0_29), .A3(n_0_28), .ZN(n_0_27));
   NOR2_X1 i_0_33 (.A1(M[17]), .A2(M[16]), .ZN(n_0_28));
   NOR2_X1 i_0_34 (.A1(M[19]), .A2(M[18]), .ZN(n_0_29));
   NOR4_X1 i_0_35 (.A1(M[23]), .A2(M[22]), .A3(M[21]), .A4(M[20]), .ZN(n_0_30));
   NOR4_X1 i_0_36 (.A1(M[11]), .A2(M[10]), .A3(M[9]), .A4(M[8]), .ZN(n_0_31));
   INV_X1 i_0_37 (.A(M[1]), .ZN(n_0_32));
   INV_X1 i_0_38 (.A(M[7]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(M[10]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(M[13]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(M[14]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(M[17]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(M[19]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(M[22]), .ZN(n_0_39));
endmodule

module datapath__0_26(A, p_0, M_temp);
   input [24:0]A;
   output [24:0]p_0;
   input [24:0]M_temp;

   INV_X1 i_0 (.A(A[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(M_temp[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(M_temp[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(A[1]), .B(M_temp[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(A[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(M_temp[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(A[2]), .B(M_temp[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(M_temp[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(A[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(A[3]), .B(M_temp[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(A[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(M_temp[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(A[4]), .B(M_temp[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(M_temp[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(A[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(A[5]), .B(M_temp[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(A[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(M_temp[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(A[6]), .B(M_temp[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(M_temp[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(A[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(A[7]), .B(M_temp[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(A[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(M_temp[7]), .ZN(n_23));
   XOR2_X1 i_32 (.A(A[8]), .B(M_temp[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_0[8]));
   INV_X1 i_34 (.A(M_temp[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(A[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(A[9]), .B(M_temp[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_0[9]));
   INV_X1 i_38 (.A(A[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(M_temp[9]), .ZN(n_29));
   XOR2_X1 i_40 (.A(A[10]), .B(M_temp[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_0[10]));
   INV_X1 i_42 (.A(M_temp[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(A[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(A[11]), .B(M_temp[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_0[11]));
   INV_X1 i_46 (.A(A[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(M_temp[11]), .ZN(n_35));
   XOR2_X1 i_48 (.A(A[12]), .B(M_temp[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_0[12]));
   INV_X1 i_50 (.A(M_temp[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(A[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(A[13]), .B(M_temp[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_0[13]));
   INV_X1 i_54 (.A(A[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(M_temp[13]), .ZN(n_41));
   XOR2_X1 i_56 (.A(A[14]), .B(M_temp[14]), .Z(n_42));
   XNOR2_X1 i_57 (.A(n_41), .B(n_42), .ZN(p_0[14]));
   INV_X1 i_58 (.A(M_temp[14]), .ZN(n_43));
   OAI22_X1 i_59 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(A[14]), .ZN(n_44));
   XNOR2_X1 i_60 (.A(A[15]), .B(M_temp[15]), .ZN(n_45));
   XNOR2_X1 i_61 (.A(n_44), .B(n_45), .ZN(p_0[15]));
   INV_X1 i_62 (.A(A[15]), .ZN(n_46));
   AOI22_X1 i_63 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(M_temp[15]), .ZN(n_47));
   XOR2_X1 i_64 (.A(A[16]), .B(M_temp[16]), .Z(n_48));
   XNOR2_X1 i_65 (.A(n_47), .B(n_48), .ZN(p_0[16]));
   INV_X1 i_66 (.A(M_temp[16]), .ZN(n_49));
   OAI22_X1 i_67 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(A[16]), .ZN(n_50));
   XNOR2_X1 i_68 (.A(A[17]), .B(M_temp[17]), .ZN(n_51));
   XNOR2_X1 i_69 (.A(n_50), .B(n_51), .ZN(p_0[17]));
   INV_X1 i_70 (.A(A[17]), .ZN(n_52));
   AOI22_X1 i_71 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(M_temp[17]), .ZN(n_53));
   XOR2_X1 i_72 (.A(A[18]), .B(M_temp[18]), .Z(n_54));
   XNOR2_X1 i_73 (.A(n_53), .B(n_54), .ZN(p_0[18]));
   INV_X1 i_74 (.A(M_temp[18]), .ZN(n_55));
   OAI22_X1 i_75 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(A[18]), .ZN(n_56));
   XNOR2_X1 i_76 (.A(A[19]), .B(M_temp[19]), .ZN(n_57));
   XNOR2_X1 i_77 (.A(n_56), .B(n_57), .ZN(p_0[19]));
   INV_X1 i_78 (.A(A[19]), .ZN(n_58));
   AOI22_X1 i_79 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(M_temp[19]), .ZN(n_59));
   XOR2_X1 i_80 (.A(A[20]), .B(M_temp[20]), .Z(n_60));
   XNOR2_X1 i_81 (.A(n_59), .B(n_60), .ZN(p_0[20]));
   INV_X1 i_82 (.A(M_temp[20]), .ZN(n_61));
   OAI22_X1 i_83 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(A[20]), .ZN(n_62));
   XNOR2_X1 i_84 (.A(A[21]), .B(M_temp[21]), .ZN(n_63));
   XNOR2_X1 i_85 (.A(n_62), .B(n_63), .ZN(p_0[21]));
   INV_X1 i_86 (.A(A[21]), .ZN(n_64));
   AOI22_X1 i_87 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(M_temp[21]), .ZN(n_65));
   XOR2_X1 i_88 (.A(A[22]), .B(M_temp[22]), .Z(n_66));
   XNOR2_X1 i_89 (.A(n_65), .B(n_66), .ZN(p_0[22]));
   INV_X1 i_90 (.A(M_temp[22]), .ZN(n_67));
   OAI22_X1 i_91 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(A[22]), .ZN(n_68));
   XNOR2_X1 i_92 (.A(A[23]), .B(M_temp[23]), .ZN(n_69));
   XNOR2_X1 i_93 (.A(n_68), .B(n_69), .ZN(p_0[23]));
   INV_X1 i_94 (.A(A[23]), .ZN(n_70));
   AOI22_X1 i_95 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(M_temp[23]), .ZN(n_71));
   XNOR2_X1 i_96 (.A(n_71), .B(A[24]), .ZN(p_0[24]));
endmodule

module datapath__0_27(M_temp, A, A0);
   input [24:0]M_temp;
   input [24:0]A;
   output [24:0]A0;

   HA_X1 i_0 (.A(M_temp[0]), .B(A[0]), .CO(n_0), .S(A0[0]));
   FA_X1 i_1 (.A(M_temp[1]), .B(A[1]), .CI(n_0), .CO(n_1), .S(A0[1]));
   FA_X1 i_2 (.A(M_temp[2]), .B(A[2]), .CI(n_1), .CO(n_2), .S(A0[2]));
   FA_X1 i_3 (.A(M_temp[3]), .B(A[3]), .CI(n_2), .CO(n_3), .S(A0[3]));
   FA_X1 i_4 (.A(M_temp[4]), .B(A[4]), .CI(n_3), .CO(n_4), .S(A0[4]));
   FA_X1 i_5 (.A(M_temp[5]), .B(A[5]), .CI(n_4), .CO(n_5), .S(A0[5]));
   FA_X1 i_6 (.A(M_temp[6]), .B(A[6]), .CI(n_5), .CO(n_6), .S(A0[6]));
   FA_X1 i_7 (.A(M_temp[7]), .B(A[7]), .CI(n_6), .CO(n_7), .S(A0[7]));
   FA_X1 i_8 (.A(M_temp[8]), .B(A[8]), .CI(n_7), .CO(n_8), .S(A0[8]));
   FA_X1 i_9 (.A(M_temp[9]), .B(A[9]), .CI(n_8), .CO(n_9), .S(A0[9]));
   FA_X1 i_10 (.A(M_temp[10]), .B(A[10]), .CI(n_9), .CO(n_10), .S(A0[10]));
   FA_X1 i_11 (.A(M_temp[11]), .B(A[11]), .CI(n_10), .CO(n_11), .S(A0[11]));
   FA_X1 i_12 (.A(M_temp[12]), .B(A[12]), .CI(n_11), .CO(n_12), .S(A0[12]));
   FA_X1 i_13 (.A(M_temp[13]), .B(A[13]), .CI(n_12), .CO(n_13), .S(A0[13]));
   FA_X1 i_14 (.A(M_temp[14]), .B(A[14]), .CI(n_13), .CO(n_14), .S(A0[14]));
   FA_X1 i_15 (.A(M_temp[15]), .B(A[15]), .CI(n_14), .CO(n_15), .S(A0[15]));
   FA_X1 i_16 (.A(M_temp[16]), .B(A[16]), .CI(n_15), .CO(n_16), .S(A0[16]));
   FA_X1 i_17 (.A(M_temp[17]), .B(A[17]), .CI(n_16), .CO(n_17), .S(A0[17]));
   FA_X1 i_18 (.A(M_temp[18]), .B(A[18]), .CI(n_17), .CO(n_18), .S(A0[18]));
   FA_X1 i_19 (.A(M_temp[19]), .B(A[19]), .CI(n_18), .CO(n_19), .S(A0[19]));
   FA_X1 i_20 (.A(M_temp[20]), .B(A[20]), .CI(n_19), .CO(n_20), .S(A0[20]));
   FA_X1 i_21 (.A(M_temp[21]), .B(A[21]), .CI(n_20), .CO(n_21), .S(A0[21]));
   FA_X1 i_22 (.A(M_temp[22]), .B(A[22]), .CI(n_21), .CO(n_22), .S(A0[22]));
   FA_X1 i_23 (.A(M_temp[23]), .B(A[23]), .CI(n_22), .CO(n_23), .S(A0[23]));
   XOR2_X1 i_24 (.A(A[24]), .B(n_23), .Z(A0[24]));
endmodule

module both_f(i_clk, i_load, i_rst, M, Q, P);
   input i_clk;
   input i_load;
   input i_rst;
   input [24:0]M;
   input [24:0]Q;
   output [47:0]P;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire [24:0]Q_temp;
   wire Q_minus_one;
   wire [4:0]Count;
   wire [24:0]M_temp;
   wire [24:0]A;

   datapath__0_26 i_6 (.A({A[24], A[23], P[47], P[46], P[45], P[44], P[43], 
      P[42], P[41], P[40], P[39], P[38], P[37], P[36], P[35], P[34], P[33], 
      P[32], P[31], P[30], P[29], P[28], P[27], P[26], P[25]}), .p_0({n_24, n_23, 
      n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
      n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .M_temp({uc_0, 
      M_temp[23], M_temp[22], M_temp[21], M_temp[20], M_temp[19], M_temp[18], 
      M_temp[17], M_temp[16], M_temp[15], M_temp[14], M_temp[13], M_temp[12], 
      M_temp[11], M_temp[10], M_temp[9], M_temp[8], M_temp[7], M_temp[6], 
      M_temp[5], M_temp[4], M_temp[3], M_temp[2], M_temp[1], M_temp[0]}));
   datapath__0_27 i_7 (.M_temp({uc_1, M_temp[23], M_temp[22], M_temp[21], 
      M_temp[20], M_temp[19], M_temp[18], M_temp[17], M_temp[16], M_temp[15], 
      M_temp[14], M_temp[13], M_temp[12], M_temp[11], M_temp[10], M_temp[9], 
      M_temp[8], M_temp[7], M_temp[6], M_temp[5], M_temp[4], M_temp[3], 
      M_temp[2], M_temp[1], M_temp[0]}), .A({A[24], A[23], P[47], P[46], P[45], 
      P[44], P[43], P[42], P[41], P[40], P[39], P[38], P[37], P[36], P[35], 
      P[34], P[33], P[32], P[31], P[30], P[29], P[28], P[27], P[26], P[25]}), 
      .A0({n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, 
      n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, 
      n_26, n_25}));
   AND2_X1 i_0_0 (.A1(n_0_92), .A2(M[0]), .ZN(n_50));
   AND2_X1 i_0_1 (.A1(n_0_92), .A2(M[1]), .ZN(n_51));
   AND2_X1 i_0_2 (.A1(n_0_92), .A2(M[2]), .ZN(n_52));
   AND2_X1 i_0_3 (.A1(n_0_92), .A2(M[3]), .ZN(n_53));
   AND2_X1 i_0_4 (.A1(n_0_92), .A2(M[4]), .ZN(n_54));
   AND2_X1 i_0_5 (.A1(n_0_92), .A2(M[5]), .ZN(n_55));
   AND2_X1 i_0_6 (.A1(n_0_92), .A2(M[6]), .ZN(n_56));
   AND2_X1 i_0_7 (.A1(n_0_92), .A2(M[7]), .ZN(n_57));
   AND2_X1 i_0_8 (.A1(n_0_92), .A2(M[8]), .ZN(n_58));
   AND2_X1 i_0_9 (.A1(n_0_92), .A2(M[9]), .ZN(n_59));
   AND2_X1 i_0_10 (.A1(n_0_92), .A2(M[10]), .ZN(n_60));
   AND2_X1 i_0_11 (.A1(n_0_92), .A2(M[11]), .ZN(n_61));
   AND2_X1 i_0_12 (.A1(n_0_92), .A2(M[12]), .ZN(n_62));
   AND2_X1 i_0_13 (.A1(n_0_92), .A2(M[13]), .ZN(n_63));
   AND2_X1 i_0_14 (.A1(n_0_92), .A2(M[14]), .ZN(n_64));
   AND2_X1 i_0_15 (.A1(n_0_92), .A2(M[15]), .ZN(n_65));
   AND2_X1 i_0_16 (.A1(n_0_92), .A2(M[16]), .ZN(n_66));
   AND2_X1 i_0_17 (.A1(n_0_92), .A2(M[17]), .ZN(n_67));
   AND2_X1 i_0_18 (.A1(n_0_92), .A2(M[18]), .ZN(n_68));
   AND2_X1 i_0_19 (.A1(n_0_92), .A2(M[19]), .ZN(n_69));
   AND2_X1 i_0_20 (.A1(n_0_92), .A2(M[20]), .ZN(n_70));
   AND2_X1 i_0_21 (.A1(n_0_92), .A2(M[21]), .ZN(n_71));
   AND2_X1 i_0_22 (.A1(n_0_92), .A2(M[22]), .ZN(n_72));
   AND2_X1 i_0_23 (.A1(n_0_92), .A2(M[23]), .ZN(n_73));
   NAND2_X1 i_0_24 (.A1(n_0_92), .A2(Count[0]), .ZN(n_74));
   NOR2_X1 i_0_25 (.A1(i_rst), .A2(n_0_0), .ZN(n_75));
   XOR2_X1 i_0_26 (.A(Count[1]), .B(Count[0]), .Z(n_0_0));
   AOI21_X1 i_0_27 (.A(i_rst), .B1(n_0_91), .B2(n_0_1), .ZN(n_76));
   OAI21_X1 i_0_28 (.A(Count[2]), .B1(Count[1]), .B2(Count[0]), .ZN(n_0_1));
   NAND2_X1 i_0_29 (.A1(n_0_90), .A2(n_0_2), .ZN(n_77));
   AOI21_X1 i_0_30 (.A(i_rst), .B1(n_0_91), .B2(Count[3]), .ZN(n_0_2));
   OAI21_X1 i_0_31 (.A(n_0_3), .B1(n_0_90), .B2(Count[4]), .ZN(n_78));
   AOI21_X1 i_0_32 (.A(i_rst), .B1(n_0_90), .B2(Count[4]), .ZN(n_0_3));
   NAND2_X1 i_0_33 (.A1(n_0_6), .A2(n_0_4), .ZN(n_79));
   AOI22_X1 i_0_34 (.A1(A[23]), .A2(n_0_84), .B1(n_0_82), .B2(A[24]), .ZN(n_0_4));
   NAND2_X1 i_0_35 (.A1(n_0_6), .A2(n_0_5), .ZN(n_80));
   NAND3_X1 i_0_36 (.A1(n_0_86), .A2(A[24]), .A3(n_0_92), .ZN(n_0_5));
   AOI22_X1 i_0_37 (.A1(n_24), .A2(n_0_85), .B1(n_0_81), .B2(n_49), .ZN(n_0_6));
   INV_X1 i_0_38 (.A(n_0_7), .ZN(n_81));
   AOI222_X1 i_0_39 (.A1(Q_temp[1]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[0]), 
      .C1(n_0_31), .C2(Q[0]), .ZN(n_0_7));
   INV_X1 i_0_40 (.A(n_0_8), .ZN(n_82));
   AOI222_X1 i_0_41 (.A1(Q_temp[2]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[1]), 
      .C1(n_0_31), .C2(Q[1]), .ZN(n_0_8));
   INV_X1 i_0_42 (.A(n_0_9), .ZN(n_83));
   AOI222_X1 i_0_43 (.A1(Q_temp[3]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[2]), 
      .C1(n_0_31), .C2(Q[2]), .ZN(n_0_9));
   INV_X1 i_0_44 (.A(n_0_10), .ZN(n_84));
   AOI222_X1 i_0_45 (.A1(Q_temp[4]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[3]), 
      .C1(n_0_31), .C2(Q[3]), .ZN(n_0_10));
   INV_X1 i_0_46 (.A(n_0_11), .ZN(n_85));
   AOI222_X1 i_0_47 (.A1(Q_temp[5]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[4]), 
      .C1(n_0_31), .C2(Q[4]), .ZN(n_0_11));
   INV_X1 i_0_48 (.A(n_0_12), .ZN(n_86));
   AOI222_X1 i_0_49 (.A1(Q_temp[6]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[5]), 
      .C1(n_0_31), .C2(Q[5]), .ZN(n_0_12));
   INV_X1 i_0_50 (.A(n_0_13), .ZN(n_87));
   AOI222_X1 i_0_51 (.A1(Q_temp[7]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[6]), 
      .C1(n_0_31), .C2(Q[6]), .ZN(n_0_13));
   INV_X1 i_0_52 (.A(n_0_14), .ZN(n_88));
   AOI222_X1 i_0_53 (.A1(Q_temp[8]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[7]), 
      .C1(n_0_31), .C2(Q[7]), .ZN(n_0_14));
   INV_X1 i_0_54 (.A(n_0_15), .ZN(n_89));
   AOI222_X1 i_0_55 (.A1(Q_temp[9]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[8]), 
      .C1(n_0_31), .C2(Q[8]), .ZN(n_0_15));
   INV_X1 i_0_56 (.A(n_0_16), .ZN(n_90));
   AOI222_X1 i_0_57 (.A1(Q_temp[10]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[9]), 
      .C1(n_0_31), .C2(Q[9]), .ZN(n_0_16));
   INV_X1 i_0_58 (.A(n_0_17), .ZN(n_91));
   AOI222_X1 i_0_59 (.A1(Q_temp[11]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[10]), 
      .C1(n_0_31), .C2(Q[10]), .ZN(n_0_17));
   INV_X1 i_0_60 (.A(n_0_18), .ZN(n_92));
   AOI222_X1 i_0_61 (.A1(Q_temp[12]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[11]), 
      .C1(n_0_31), .C2(Q[11]), .ZN(n_0_18));
   INV_X1 i_0_62 (.A(n_0_19), .ZN(n_93));
   AOI222_X1 i_0_63 (.A1(Q_temp[13]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[12]), 
      .C1(n_0_31), .C2(Q[12]), .ZN(n_0_19));
   INV_X1 i_0_64 (.A(n_0_20), .ZN(n_94));
   AOI222_X1 i_0_65 (.A1(Q_temp[14]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[13]), 
      .C1(n_0_31), .C2(Q[13]), .ZN(n_0_20));
   INV_X1 i_0_66 (.A(n_0_21), .ZN(n_95));
   AOI222_X1 i_0_67 (.A1(Q_temp[15]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[14]), 
      .C1(n_0_31), .C2(Q[14]), .ZN(n_0_21));
   INV_X1 i_0_68 (.A(n_0_22), .ZN(n_96));
   AOI222_X1 i_0_69 (.A1(Q_temp[16]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[15]), 
      .C1(n_0_31), .C2(Q[15]), .ZN(n_0_22));
   INV_X1 i_0_70 (.A(n_0_23), .ZN(n_97));
   AOI222_X1 i_0_71 (.A1(Q_temp[17]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[16]), 
      .C1(n_0_31), .C2(Q[16]), .ZN(n_0_23));
   INV_X1 i_0_72 (.A(n_0_24), .ZN(n_98));
   AOI222_X1 i_0_73 (.A1(Q_temp[18]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[17]), 
      .C1(n_0_31), .C2(Q[17]), .ZN(n_0_24));
   INV_X1 i_0_74 (.A(n_0_25), .ZN(n_99));
   AOI222_X1 i_0_75 (.A1(Q_temp[19]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[18]), 
      .C1(n_0_31), .C2(Q[18]), .ZN(n_0_25));
   INV_X1 i_0_76 (.A(n_0_26), .ZN(n_100));
   AOI222_X1 i_0_77 (.A1(Q_temp[20]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[19]), 
      .C1(n_0_31), .C2(Q[19]), .ZN(n_0_26));
   INV_X1 i_0_78 (.A(n_0_27), .ZN(n_101));
   AOI222_X1 i_0_79 (.A1(Q_temp[21]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[20]), 
      .C1(n_0_31), .C2(Q[20]), .ZN(n_0_27));
   INV_X1 i_0_80 (.A(n_0_28), .ZN(n_102));
   AOI222_X1 i_0_81 (.A1(Q_temp[22]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[21]), 
      .C1(n_0_31), .C2(Q[21]), .ZN(n_0_28));
   INV_X1 i_0_82 (.A(n_0_29), .ZN(n_103));
   AOI222_X1 i_0_83 (.A1(P[23]), .A2(n_0_83), .B1(n_0_34), .B2(Q_temp[22]), 
      .C1(n_0_31), .C2(Q[22]), .ZN(n_0_29));
   INV_X1 i_0_84 (.A(n_0_30), .ZN(n_104));
   AOI222_X1 i_0_85 (.A1(P[24]), .A2(n_0_83), .B1(n_0_34), .B2(P[23]), .C1(
      n_0_31), .C2(Q[23]), .ZN(n_0_30));
   AND2_X1 i_0_86 (.A1(n_0_92), .A2(i_load), .ZN(n_0_31));
   NAND2_X1 i_0_87 (.A1(n_0_33), .A2(n_0_32), .ZN(n_105));
   AOI22_X1 i_0_88 (.A1(n_0), .A2(n_0_85), .B1(n_0_34), .B2(P[24]), .ZN(n_0_32));
   AOI22_X1 i_0_89 (.A1(P[25]), .A2(n_0_82), .B1(n_0_81), .B2(n_25), .ZN(n_0_33));
   NOR3_X1 i_0_90 (.A1(n_0_90), .A2(n_129), .A3(Count[4]), .ZN(n_0_34));
   NAND2_X1 i_0_91 (.A1(n_0_36), .A2(n_0_35), .ZN(n_106));
   AOI22_X1 i_0_92 (.A1(n_1), .A2(n_0_85), .B1(n_0_81), .B2(n_26), .ZN(n_0_35));
   AOI22_X1 i_0_93 (.A1(P[25]), .A2(n_0_84), .B1(n_0_82), .B2(P[26]), .ZN(n_0_36));
   NAND2_X1 i_0_94 (.A1(n_0_38), .A2(n_0_37), .ZN(n_107));
   AOI22_X1 i_0_95 (.A1(n_2), .A2(n_0_85), .B1(n_0_81), .B2(n_27), .ZN(n_0_37));
   AOI22_X1 i_0_96 (.A1(P[26]), .A2(n_0_84), .B1(n_0_82), .B2(P[27]), .ZN(n_0_38));
   NAND2_X1 i_0_97 (.A1(n_0_40), .A2(n_0_39), .ZN(n_108));
   AOI22_X1 i_0_98 (.A1(n_3), .A2(n_0_85), .B1(n_0_81), .B2(n_28), .ZN(n_0_39));
   AOI22_X1 i_0_99 (.A1(P[27]), .A2(n_0_84), .B1(n_0_82), .B2(P[28]), .ZN(n_0_40));
   NAND2_X1 i_0_100 (.A1(n_0_42), .A2(n_0_41), .ZN(n_109));
   AOI22_X1 i_0_101 (.A1(n_4), .A2(n_0_85), .B1(n_0_81), .B2(n_29), .ZN(n_0_41));
   AOI22_X1 i_0_102 (.A1(P[28]), .A2(n_0_84), .B1(n_0_82), .B2(P[29]), .ZN(
      n_0_42));
   NAND2_X1 i_0_103 (.A1(n_0_44), .A2(n_0_43), .ZN(n_110));
   AOI22_X1 i_0_104 (.A1(n_5), .A2(n_0_85), .B1(n_0_81), .B2(n_30), .ZN(n_0_43));
   AOI22_X1 i_0_105 (.A1(P[29]), .A2(n_0_84), .B1(n_0_82), .B2(P[30]), .ZN(
      n_0_44));
   NAND2_X1 i_0_106 (.A1(n_0_46), .A2(n_0_45), .ZN(n_111));
   AOI22_X1 i_0_107 (.A1(n_6), .A2(n_0_85), .B1(n_0_81), .B2(n_31), .ZN(n_0_45));
   AOI22_X1 i_0_108 (.A1(P[30]), .A2(n_0_84), .B1(n_0_82), .B2(P[31]), .ZN(
      n_0_46));
   NAND2_X1 i_0_109 (.A1(n_0_48), .A2(n_0_47), .ZN(n_112));
   AOI22_X1 i_0_110 (.A1(n_7), .A2(n_0_85), .B1(n_0_81), .B2(n_32), .ZN(n_0_47));
   AOI22_X1 i_0_111 (.A1(P[31]), .A2(n_0_84), .B1(n_0_82), .B2(P[32]), .ZN(
      n_0_48));
   NAND2_X1 i_0_112 (.A1(n_0_50), .A2(n_0_49), .ZN(n_113));
   AOI22_X1 i_0_113 (.A1(n_8), .A2(n_0_85), .B1(n_0_81), .B2(n_33), .ZN(n_0_49));
   AOI22_X1 i_0_114 (.A1(P[32]), .A2(n_0_84), .B1(n_0_82), .B2(P[33]), .ZN(
      n_0_50));
   NAND2_X1 i_0_115 (.A1(n_0_52), .A2(n_0_51), .ZN(n_114));
   AOI22_X1 i_0_116 (.A1(n_9), .A2(n_0_85), .B1(n_0_81), .B2(n_34), .ZN(n_0_51));
   AOI22_X1 i_0_117 (.A1(P[33]), .A2(n_0_84), .B1(n_0_82), .B2(P[34]), .ZN(
      n_0_52));
   NAND2_X1 i_0_118 (.A1(n_0_54), .A2(n_0_53), .ZN(n_115));
   AOI22_X1 i_0_119 (.A1(n_10), .A2(n_0_85), .B1(n_0_81), .B2(n_35), .ZN(n_0_53));
   AOI22_X1 i_0_120 (.A1(P[34]), .A2(n_0_84), .B1(n_0_82), .B2(P[35]), .ZN(
      n_0_54));
   NAND2_X1 i_0_121 (.A1(n_0_56), .A2(n_0_55), .ZN(n_116));
   AOI22_X1 i_0_122 (.A1(n_11), .A2(n_0_85), .B1(n_0_81), .B2(n_36), .ZN(n_0_55));
   AOI22_X1 i_0_123 (.A1(P[35]), .A2(n_0_84), .B1(n_0_82), .B2(P[36]), .ZN(
      n_0_56));
   NAND2_X1 i_0_124 (.A1(n_0_58), .A2(n_0_57), .ZN(n_117));
   AOI22_X1 i_0_125 (.A1(n_12), .A2(n_0_85), .B1(n_0_81), .B2(n_37), .ZN(n_0_57));
   AOI22_X1 i_0_126 (.A1(P[36]), .A2(n_0_84), .B1(n_0_82), .B2(P[37]), .ZN(
      n_0_58));
   NAND2_X1 i_0_127 (.A1(n_0_60), .A2(n_0_59), .ZN(n_118));
   AOI22_X1 i_0_128 (.A1(n_13), .A2(n_0_85), .B1(n_0_81), .B2(n_38), .ZN(n_0_59));
   AOI22_X1 i_0_129 (.A1(P[37]), .A2(n_0_84), .B1(n_0_82), .B2(P[38]), .ZN(
      n_0_60));
   NAND2_X1 i_0_130 (.A1(n_0_62), .A2(n_0_61), .ZN(n_119));
   AOI22_X1 i_0_131 (.A1(n_14), .A2(n_0_85), .B1(n_0_81), .B2(n_39), .ZN(n_0_61));
   AOI22_X1 i_0_132 (.A1(P[38]), .A2(n_0_84), .B1(n_0_82), .B2(P[39]), .ZN(
      n_0_62));
   NAND2_X1 i_0_133 (.A1(n_0_64), .A2(n_0_63), .ZN(n_120));
   AOI22_X1 i_0_134 (.A1(n_15), .A2(n_0_85), .B1(n_0_81), .B2(n_40), .ZN(n_0_63));
   AOI22_X1 i_0_135 (.A1(P[39]), .A2(n_0_84), .B1(n_0_82), .B2(P[40]), .ZN(
      n_0_64));
   NAND2_X1 i_0_136 (.A1(n_0_66), .A2(n_0_65), .ZN(n_121));
   AOI22_X1 i_0_137 (.A1(n_16), .A2(n_0_85), .B1(n_0_81), .B2(n_41), .ZN(n_0_65));
   AOI22_X1 i_0_138 (.A1(P[40]), .A2(n_0_84), .B1(n_0_82), .B2(P[41]), .ZN(
      n_0_66));
   NAND2_X1 i_0_139 (.A1(n_0_68), .A2(n_0_67), .ZN(n_122));
   AOI22_X1 i_0_140 (.A1(n_17), .A2(n_0_85), .B1(n_0_81), .B2(n_42), .ZN(n_0_67));
   AOI22_X1 i_0_141 (.A1(P[41]), .A2(n_0_84), .B1(n_0_82), .B2(P[42]), .ZN(
      n_0_68));
   NAND2_X1 i_0_142 (.A1(n_0_70), .A2(n_0_69), .ZN(n_123));
   AOI22_X1 i_0_143 (.A1(n_18), .A2(n_0_85), .B1(n_0_81), .B2(n_43), .ZN(n_0_69));
   AOI22_X1 i_0_144 (.A1(P[42]), .A2(n_0_84), .B1(n_0_82), .B2(P[43]), .ZN(
      n_0_70));
   NAND2_X1 i_0_145 (.A1(n_0_72), .A2(n_0_71), .ZN(n_124));
   AOI22_X1 i_0_146 (.A1(n_19), .A2(n_0_85), .B1(n_0_81), .B2(n_44), .ZN(n_0_71));
   AOI22_X1 i_0_147 (.A1(P[43]), .A2(n_0_84), .B1(n_0_82), .B2(P[44]), .ZN(
      n_0_72));
   NAND2_X1 i_0_148 (.A1(n_0_74), .A2(n_0_73), .ZN(n_125));
   AOI22_X1 i_0_149 (.A1(n_20), .A2(n_0_85), .B1(n_0_81), .B2(n_45), .ZN(n_0_73));
   AOI22_X1 i_0_150 (.A1(P[44]), .A2(n_0_84), .B1(n_0_82), .B2(P[45]), .ZN(
      n_0_74));
   NAND2_X1 i_0_151 (.A1(n_0_76), .A2(n_0_75), .ZN(n_126));
   AOI22_X1 i_0_152 (.A1(n_21), .A2(n_0_85), .B1(n_0_81), .B2(n_46), .ZN(n_0_75));
   AOI22_X1 i_0_153 (.A1(P[45]), .A2(n_0_84), .B1(n_0_82), .B2(P[46]), .ZN(
      n_0_76));
   NAND2_X1 i_0_154 (.A1(n_0_78), .A2(n_0_77), .ZN(n_127));
   AOI22_X1 i_0_155 (.A1(n_22), .A2(n_0_85), .B1(n_0_81), .B2(n_47), .ZN(n_0_77));
   AOI22_X1 i_0_156 (.A1(P[46]), .A2(n_0_84), .B1(n_0_82), .B2(P[47]), .ZN(
      n_0_78));
   NAND2_X1 i_0_157 (.A1(n_0_80), .A2(n_0_79), .ZN(n_128));
   AOI22_X1 i_0_158 (.A1(n_23), .A2(n_0_85), .B1(n_0_81), .B2(n_48), .ZN(n_0_79));
   AOI22_X1 i_0_159 (.A1(P[47]), .A2(n_0_84), .B1(n_0_82), .B2(A[23]), .ZN(
      n_0_80));
   AND3_X1 i_0_160 (.A1(Q_minus_one), .A2(n_0_83), .A3(n_0_93), .ZN(n_0_81));
   NOR3_X1 i_0_161 (.A1(n_0_89), .A2(n_0_87), .A3(n_129), .ZN(n_0_82));
   NOR2_X1 i_0_162 (.A1(n_0_89), .A2(n_129), .ZN(n_0_83));
   OR2_X1 i_0_163 (.A1(i_rst), .A2(i_load), .ZN(n_129));
   INV_X1 i_0_164 (.A(n_0_84), .ZN(n_130));
   NOR2_X1 i_0_165 (.A1(i_rst), .A2(n_0_88), .ZN(n_0_84));
   NOR3_X1 i_0_166 (.A1(n_0_93), .A2(n_0_86), .A3(i_rst), .ZN(n_0_85));
   NAND2_X1 i_0_167 (.A1(n_0_88), .A2(n_0_87), .ZN(n_0_86));
   XNOR2_X1 i_0_168 (.A(Q_minus_one), .B(n_0_93), .ZN(n_0_87));
   NOR2_X1 i_0_169 (.A1(i_load), .A2(n_0_89), .ZN(n_0_88));
   NOR2_X1 i_0_170 (.A1(n_0_90), .A2(Count[4]), .ZN(n_0_89));
   OR2_X1 i_0_171 (.A1(n_0_91), .A2(Count[3]), .ZN(n_0_90));
   OR3_X1 i_0_172 (.A1(Count[2]), .A2(Count[1]), .A3(Count[0]), .ZN(n_0_91));
   NOR2_X1 i_0_173 (.A1(n_0_93), .A2(i_rst), .ZN(n_131));
   INV_X1 i_0_174 (.A(i_rst), .ZN(n_0_92));
   INV_X1 i_0_175 (.A(Q_temp[0]), .ZN(n_0_93));
   DFF_X1 \Q_temp_reg[22]  (.D(n_103), .CK(i_clk), .Q(Q_temp[22]), .QN());
   DFF_X1 \Q_temp_reg[21]  (.D(n_102), .CK(i_clk), .Q(Q_temp[21]), .QN());
   DFF_X1 \Q_temp_reg[20]  (.D(n_101), .CK(i_clk), .Q(Q_temp[20]), .QN());
   DFF_X1 \Q_temp_reg[19]  (.D(n_100), .CK(i_clk), .Q(Q_temp[19]), .QN());
   DFF_X1 \Q_temp_reg[18]  (.D(n_99), .CK(i_clk), .Q(Q_temp[18]), .QN());
   DFF_X1 \Q_temp_reg[17]  (.D(n_98), .CK(i_clk), .Q(Q_temp[17]), .QN());
   DFF_X1 \Q_temp_reg[16]  (.D(n_97), .CK(i_clk), .Q(Q_temp[16]), .QN());
   DFF_X1 \Q_temp_reg[15]  (.D(n_96), .CK(i_clk), .Q(Q_temp[15]), .QN());
   DFF_X1 \Q_temp_reg[14]  (.D(n_95), .CK(i_clk), .Q(Q_temp[14]), .QN());
   DFF_X1 \Q_temp_reg[13]  (.D(n_94), .CK(i_clk), .Q(Q_temp[13]), .QN());
   DFF_X1 \Q_temp_reg[12]  (.D(n_93), .CK(i_clk), .Q(Q_temp[12]), .QN());
   DFF_X1 \Q_temp_reg[11]  (.D(n_92), .CK(i_clk), .Q(Q_temp[11]), .QN());
   DFF_X1 \Q_temp_reg[10]  (.D(n_91), .CK(i_clk), .Q(Q_temp[10]), .QN());
   DFF_X1 \Q_temp_reg[9]  (.D(n_90), .CK(i_clk), .Q(Q_temp[9]), .QN());
   DFF_X1 \Q_temp_reg[8]  (.D(n_89), .CK(i_clk), .Q(Q_temp[8]), .QN());
   DFF_X1 \Q_temp_reg[7]  (.D(n_88), .CK(i_clk), .Q(Q_temp[7]), .QN());
   DFF_X1 \Q_temp_reg[6]  (.D(n_87), .CK(i_clk), .Q(Q_temp[6]), .QN());
   DFF_X1 \Q_temp_reg[5]  (.D(n_86), .CK(i_clk), .Q(Q_temp[5]), .QN());
   DFF_X1 \Q_temp_reg[4]  (.D(n_85), .CK(i_clk), .Q(Q_temp[4]), .QN());
   DFF_X1 \Q_temp_reg[3]  (.D(n_84), .CK(i_clk), .Q(Q_temp[3]), .QN());
   DFF_X1 \Q_temp_reg[2]  (.D(n_83), .CK(i_clk), .Q(Q_temp[2]), .QN());
   DFF_X1 \Q_temp_reg[1]  (.D(n_82), .CK(i_clk), .Q(Q_temp[1]), .QN());
   DFF_X1 \Q_temp_reg[0]  (.D(n_81), .CK(i_clk), .Q(Q_temp[0]), .QN());
   DFF_X1 Q_minus_one_reg (.D(n_131), .CK(n_133), .Q(Q_minus_one), .QN());
   DFF_X1 \Count_reg[4]  (.D(n_78), .CK(n_133), .Q(Count[4]), .QN());
   DFF_X1 \Count_reg[3]  (.D(n_77), .CK(n_133), .Q(Count[3]), .QN());
   DFF_X1 \Count_reg[2]  (.D(n_76), .CK(n_133), .Q(Count[2]), .QN());
   DFF_X1 \Count_reg[1]  (.D(n_75), .CK(n_133), .Q(Count[1]), .QN());
   DFF_X1 \Count_reg[0]  (.D(n_74), .CK(n_133), .Q(Count[0]), .QN());
   CLKGATETST_X1 clk_gate_M_temp_reg (.CK(i_clk), .E(n_129), .SE(1'b0), .GCK(
      n_132));
   DFF_X1 \M_temp_reg[23]  (.D(n_73), .CK(n_132), .Q(M_temp[23]), .QN());
   DFF_X1 \M_temp_reg[22]  (.D(n_72), .CK(n_132), .Q(M_temp[22]), .QN());
   DFF_X1 \M_temp_reg[21]  (.D(n_71), .CK(n_132), .Q(M_temp[21]), .QN());
   DFF_X1 \M_temp_reg[20]  (.D(n_70), .CK(n_132), .Q(M_temp[20]), .QN());
   DFF_X1 \M_temp_reg[19]  (.D(n_69), .CK(n_132), .Q(M_temp[19]), .QN());
   DFF_X1 \M_temp_reg[18]  (.D(n_68), .CK(n_132), .Q(M_temp[18]), .QN());
   DFF_X1 \M_temp_reg[17]  (.D(n_67), .CK(n_132), .Q(M_temp[17]), .QN());
   DFF_X1 \M_temp_reg[16]  (.D(n_66), .CK(n_132), .Q(M_temp[16]), .QN());
   DFF_X1 \M_temp_reg[15]  (.D(n_65), .CK(n_132), .Q(M_temp[15]), .QN());
   DFF_X1 \M_temp_reg[14]  (.D(n_64), .CK(n_132), .Q(M_temp[14]), .QN());
   DFF_X1 \M_temp_reg[13]  (.D(n_63), .CK(n_132), .Q(M_temp[13]), .QN());
   DFF_X1 \M_temp_reg[12]  (.D(n_62), .CK(n_132), .Q(M_temp[12]), .QN());
   DFF_X1 \M_temp_reg[11]  (.D(n_61), .CK(n_132), .Q(M_temp[11]), .QN());
   DFF_X1 \M_temp_reg[10]  (.D(n_60), .CK(n_132), .Q(M_temp[10]), .QN());
   DFF_X1 \M_temp_reg[9]  (.D(n_59), .CK(n_132), .Q(M_temp[9]), .QN());
   DFF_X1 \M_temp_reg[8]  (.D(n_58), .CK(n_132), .Q(M_temp[8]), .QN());
   DFF_X1 \M_temp_reg[7]  (.D(n_57), .CK(n_132), .Q(M_temp[7]), .QN());
   DFF_X1 \M_temp_reg[6]  (.D(n_56), .CK(n_132), .Q(M_temp[6]), .QN());
   DFF_X1 \M_temp_reg[5]  (.D(n_55), .CK(n_132), .Q(M_temp[5]), .QN());
   DFF_X1 \M_temp_reg[4]  (.D(n_54), .CK(n_132), .Q(M_temp[4]), .QN());
   DFF_X1 \M_temp_reg[3]  (.D(n_53), .CK(n_132), .Q(M_temp[3]), .QN());
   DFF_X1 \M_temp_reg[2]  (.D(n_52), .CK(n_132), .Q(M_temp[2]), .QN());
   DFF_X1 \M_temp_reg[1]  (.D(n_51), .CK(n_132), .Q(M_temp[1]), .QN());
   DFF_X1 \M_temp_reg[0]  (.D(n_50), .CK(n_132), .Q(M_temp[0]), .QN());
   DFF_X1 \A_reg[24]  (.D(n_80), .CK(i_clk), .Q(A[24]), .QN());
   DFF_X1 \A_reg[23]  (.D(n_79), .CK(i_clk), .Q(A[23]), .QN());
   CLKGATETST_X1 clk_gate_Q_minus_one_reg (.CK(i_clk), .E(n_130), .SE(1'b0), 
      .GCK(n_133));
   DFF_X1 \P_reg[23]  (.D(n_104), .CK(i_clk), .Q(P[23]), .QN());
   DFF_X1 \P_reg[24]  (.D(n_105), .CK(i_clk), .Q(P[24]), .QN());
   DFF_X1 \P_reg[25]  (.D(n_106), .CK(i_clk), .Q(P[25]), .QN());
   DFF_X1 \P_reg[26]  (.D(n_107), .CK(i_clk), .Q(P[26]), .QN());
   DFF_X1 \P_reg[27]  (.D(n_108), .CK(i_clk), .Q(P[27]), .QN());
   DFF_X1 \P_reg[28]  (.D(n_109), .CK(i_clk), .Q(P[28]), .QN());
   DFF_X1 \P_reg[29]  (.D(n_110), .CK(i_clk), .Q(P[29]), .QN());
   DFF_X1 \P_reg[30]  (.D(n_111), .CK(i_clk), .Q(P[30]), .QN());
   DFF_X1 \P_reg[31]  (.D(n_112), .CK(i_clk), .Q(P[31]), .QN());
   DFF_X1 \P_reg[32]  (.D(n_113), .CK(i_clk), .Q(P[32]), .QN());
   DFF_X1 \P_reg[33]  (.D(n_114), .CK(i_clk), .Q(P[33]), .QN());
   DFF_X1 \P_reg[34]  (.D(n_115), .CK(i_clk), .Q(P[34]), .QN());
   DFF_X1 \P_reg[35]  (.D(n_116), .CK(i_clk), .Q(P[35]), .QN());
   DFF_X1 \P_reg[36]  (.D(n_117), .CK(i_clk), .Q(P[36]), .QN());
   DFF_X1 \P_reg[37]  (.D(n_118), .CK(i_clk), .Q(P[37]), .QN());
   DFF_X1 \P_reg[38]  (.D(n_119), .CK(i_clk), .Q(P[38]), .QN());
   DFF_X1 \P_reg[39]  (.D(n_120), .CK(i_clk), .Q(P[39]), .QN());
   DFF_X1 \P_reg[40]  (.D(n_121), .CK(i_clk), .Q(P[40]), .QN());
   DFF_X1 \P_reg[41]  (.D(n_122), .CK(i_clk), .Q(P[41]), .QN());
   DFF_X1 \P_reg[42]  (.D(n_123), .CK(i_clk), .Q(P[42]), .QN());
   DFF_X1 \P_reg[43]  (.D(n_124), .CK(i_clk), .Q(P[43]), .QN());
   DFF_X1 \P_reg[44]  (.D(n_125), .CK(i_clk), .Q(P[44]), .QN());
   DFF_X1 \P_reg[45]  (.D(n_126), .CK(i_clk), .Q(P[45]), .QN());
   DFF_X1 \P_reg[46]  (.D(n_127), .CK(i_clk), .Q(P[46]), .QN());
   DFF_X1 \P_reg[47]  (.D(n_128), .CK(i_clk), .Q(P[47]), .QN());
endmodule

module floating(i_clk, i_rst, i_load, i_a, i_b, o_res, o_overflow, o_underflow);
   input i_clk;
   input i_rst;
   input i_load;
   input [31:0]i_a;
   input [31:0]i_b;
   output [31:0]o_res;
   output o_overflow;
   output o_underflow;

   wire enable;
   wire [2:0]outB;
   wire [2:0]outA;
   wire [31:0]special_res;
   wire [4:0]shamt;
   wire [47:0]mult_res;
   wire Sb;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire b;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire Sa;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire [8:0]E_sum;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_12;
   wire n_0_0_7;
   wire n_0_0_13;
   wire n_0_0_8;
   wire n_0_0_14;
   wire n_0_0_9;
   wire n_0_0_15;
   wire n_0_0_10;
   wire n_0_0_16;
   wire n_0_0_11;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire [7:0]Eb;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire [23:0]Na;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire [31:0]res;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_62;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_266;
   wire n_0_0_267;
   wire [23:0]Nb;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_329;
   wire n_0_0_332;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_81;
   wire n_0_0_369;
   wire n_0_65;
   wire n_0_0_371;
   wire n_0_69;
   wire n_0_0_372;
   wire n_0_85;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_63;
   wire n_0_0_381;
   wire n_0_0_383;
   wire n_0_67;
   wire n_0_0_384;
   wire n_0_83;
   wire n_0_0_385;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_391;
   wire n_0_66;
   wire n_0_0_392;
   wire n_0_82;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_86;
   wire n_0_0_397;
   wire n_0_0_399;
   wire n_0_64;
   wire n_0_0_401;
   wire n_0_0_403;
   wire n_0_0_405;
   wire n_0_68;
   wire n_0_0_406;
   wire n_0_84;
   wire n_0_0_408;
   wire n_0_0_28;
   wire n_0_0_63;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_61;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_134;
   wire n_0_0_140;
   wire n_0_0_147;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_175;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_265;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_305;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_338;
   wire n_0_0_341;
   wire n_0_0_344;
   wire n_0_0_347;
   wire n_0_0_370;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_377;
   wire n_0_0_380;
   wire n_0_0_382;
   wire n_0_0_386;
   wire n_0_0_390;
   wire n_0_0_393;
   wire n_0_0_396;
   wire n_0_0_398;
   wire n_0_0_400;
   wire n_0_0_402;
   wire n_0_0_404;
   wire n_0_0_407;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_72;
   wire n_0_0_415;
   wire n_0_73;
   wire n_0_0_416;
   wire n_0_74;
   wire n_0_0_417;
   wire n_0_76;
   wire n_0_0_418;
   wire n_0_77;
   wire n_0_0_419;
   wire n_0_78;
   wire n_0_0_420;
   wire n_0_79;
   wire n_0_0_421;
   wire n_0_80;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_75;
   wire n_0_0_426;
   wire n_0_70;
   wire n_0_0_427;
   wire n_0_71;
   wire n_0_0_428;

   n_case ncase (.A({Sa, n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, 
      n_0_37, n_0_38, n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, 
      n_0_46, n_0_47, n_0_48, n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, n_0_54, 
      n_0_55, n_0_56, n_0_57, n_0_58, n_0_59, n_0_60}), .B({Sb, n_0_0, n_0_1, 
      n_0_2, n_0_3, n_0_4, n_0_5, n_0_6, b, n_0_7, n_0_8, n_0_9, n_0_10, n_0_11, 
      n_0_12, n_0_13, n_0_14, n_0_15, n_0_16, n_0_17, n_0_18, n_0_19, n_0_20, 
      n_0_21, n_0_22, n_0_23, n_0_24, n_0_25, n_0_26, n_0_27, n_0_28, n_0_29}), 
      .S({special_res[31], special_res[23], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6, special_res[0], uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, 
      uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, 
      uc_25, uc_26, uc_27, uc_28}), .outA(outA), .outB(outB), .enable(enable));
   zero_counter zcn (.M({n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70}), .Zcount(
      shamt));
   both_f mul_unit (.i_clk(i_clk), .i_load(i_load), .i_rst(i_rst), .M({uc_29, 
      Na[23], Na[22], Na[21], Na[20], Na[19], Na[18], Na[17], Na[16], Na[15], 
      Na[14], Na[13], Na[12], Na[11], Na[10], Na[9], Na[8], Na[7], Na[6], Na[5], 
      Na[4], Na[3], Na[2], Na[1], Na[0]}), .Q({uc_30, Nb[23], Nb[22], Nb[21], 
      Nb[20], Nb[19], Nb[18], Nb[17], Nb[16], Nb[15], Nb[14], Nb[13], Nb[12], 
      Nb[11], Nb[10], Nb[9], Nb[8], Nb[7], Nb[6], Nb[5], Nb[4], Nb[3], Nb[2], 
      Nb[1], Nb[0]}), .P({mult_res[47], mult_res[46], mult_res[45], mult_res[44], 
      mult_res[43], mult_res[42], mult_res[41], mult_res[40], mult_res[39], 
      mult_res[38], mult_res[37], mult_res[36], mult_res[35], mult_res[34], 
      mult_res[33], mult_res[32], mult_res[31], mult_res[30], mult_res[29], 
      mult_res[28], mult_res[27], mult_res[26], mult_res[25], mult_res[24], 
      mult_res[23], uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, 
      uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, 
      uc_49, uc_50, uc_51, uc_52, uc_53}));
   DFF_X1 o_underflow_reg (.D(n_0_62), .CK(i_clk), .Q(o_underflow), .QN());
   DFF_X1 o_overflow_reg (.D(n_0_61), .CK(i_clk), .Q(o_overflow), .QN());
   DFF_X1 \o_res_reg[31]  (.D(res[31]), .CK(i_clk), .Q(o_res[31]), .QN());
   DFF_X1 \o_res_reg[30]  (.D(res[30]), .CK(i_clk), .Q(o_res[30]), .QN());
   DFF_X1 \o_res_reg[29]  (.D(res[29]), .CK(i_clk), .Q(o_res[29]), .QN());
   DFF_X1 \o_res_reg[28]  (.D(res[28]), .CK(i_clk), .Q(o_res[28]), .QN());
   DFF_X1 \o_res_reg[27]  (.D(res[27]), .CK(i_clk), .Q(o_res[27]), .QN());
   DFF_X1 \o_res_reg[26]  (.D(res[26]), .CK(i_clk), .Q(o_res[26]), .QN());
   DFF_X1 \o_res_reg[25]  (.D(res[25]), .CK(i_clk), .Q(o_res[25]), .QN());
   DFF_X1 \o_res_reg[24]  (.D(res[24]), .CK(i_clk), .Q(o_res[24]), .QN());
   DFF_X1 \o_res_reg[23]  (.D(res[23]), .CK(i_clk), .Q(o_res[23]), .QN());
   DFF_X1 \o_res_reg[22]  (.D(res[22]), .CK(i_clk), .Q(o_res[22]), .QN());
   DFF_X1 \o_res_reg[21]  (.D(res[21]), .CK(i_clk), .Q(o_res[21]), .QN());
   DFF_X1 \o_res_reg[20]  (.D(res[20]), .CK(i_clk), .Q(o_res[20]), .QN());
   DFF_X1 \o_res_reg[19]  (.D(res[19]), .CK(i_clk), .Q(o_res[19]), .QN());
   DFF_X1 \o_res_reg[18]  (.D(res[18]), .CK(i_clk), .Q(o_res[18]), .QN());
   DFF_X1 \o_res_reg[17]  (.D(res[17]), .CK(i_clk), .Q(o_res[17]), .QN());
   DFF_X1 \o_res_reg[16]  (.D(res[16]), .CK(i_clk), .Q(o_res[16]), .QN());
   DFF_X1 \o_res_reg[15]  (.D(res[15]), .CK(i_clk), .Q(o_res[15]), .QN());
   DFF_X1 \o_res_reg[14]  (.D(res[14]), .CK(i_clk), .Q(o_res[14]), .QN());
   DFF_X1 \o_res_reg[13]  (.D(res[13]), .CK(i_clk), .Q(o_res[13]), .QN());
   DFF_X1 \o_res_reg[12]  (.D(res[12]), .CK(i_clk), .Q(o_res[12]), .QN());
   DFF_X1 \o_res_reg[11]  (.D(res[11]), .CK(i_clk), .Q(o_res[11]), .QN());
   DFF_X1 \o_res_reg[10]  (.D(res[10]), .CK(i_clk), .Q(o_res[10]), .QN());
   DFF_X1 \o_res_reg[9]  (.D(res[9]), .CK(i_clk), .Q(o_res[9]), .QN());
   DFF_X1 \o_res_reg[8]  (.D(res[8]), .CK(i_clk), .Q(o_res[8]), .QN());
   DFF_X1 \o_res_reg[7]  (.D(res[7]), .CK(i_clk), .Q(o_res[7]), .QN());
   DFF_X1 \o_res_reg[6]  (.D(res[6]), .CK(i_clk), .Q(o_res[6]), .QN());
   DFF_X1 \o_res_reg[5]  (.D(res[5]), .CK(i_clk), .Q(o_res[5]), .QN());
   DFF_X1 \o_res_reg[4]  (.D(res[4]), .CK(i_clk), .Q(o_res[4]), .QN());
   DFF_X1 \o_res_reg[3]  (.D(res[3]), .CK(i_clk), .Q(o_res[3]), .QN());
   DFF_X1 \o_res_reg[2]  (.D(res[2]), .CK(i_clk), .Q(o_res[2]), .QN());
   DFF_X1 \o_res_reg[1]  (.D(res[1]), .CK(i_clk), .Q(o_res[1]), .QN());
   DFF_X1 \o_res_reg[0]  (.D(res[0]), .CK(i_clk), .Q(o_res[0]), .QN());
   DFF_X1 \b_reg[31]  (.D(i_b[31]), .CK(i_clk), .Q(Sb), .QN());
   DFF_X1 \b_reg[30]  (.D(i_b[30]), .CK(i_clk), .Q(n_0_0), .QN());
   DFF_X1 \b_reg[29]  (.D(i_b[29]), .CK(i_clk), .Q(n_0_1), .QN());
   DFF_X1 \b_reg[28]  (.D(i_b[28]), .CK(i_clk), .Q(n_0_2), .QN());
   DFF_X1 \b_reg[27]  (.D(i_b[27]), .CK(i_clk), .Q(n_0_3), .QN());
   DFF_X1 \b_reg[26]  (.D(i_b[26]), .CK(i_clk), .Q(n_0_4), .QN());
   DFF_X1 \b_reg[25]  (.D(i_b[25]), .CK(i_clk), .Q(n_0_5), .QN());
   DFF_X1 \b_reg[24]  (.D(i_b[24]), .CK(i_clk), .Q(n_0_6), .QN());
   DFF_X1 \b_reg[23]  (.D(i_b[23]), .CK(i_clk), .Q(b), .QN());
   DFF_X1 \b_reg[22]  (.D(i_b[22]), .CK(i_clk), .Q(n_0_7), .QN());
   DFF_X1 \b_reg[21]  (.D(i_b[21]), .CK(i_clk), .Q(n_0_8), .QN());
   DFF_X1 \b_reg[20]  (.D(i_b[20]), .CK(i_clk), .Q(n_0_9), .QN());
   DFF_X1 \b_reg[19]  (.D(i_b[19]), .CK(i_clk), .Q(n_0_10), .QN());
   DFF_X1 \b_reg[18]  (.D(i_b[18]), .CK(i_clk), .Q(n_0_11), .QN());
   DFF_X1 \b_reg[17]  (.D(i_b[17]), .CK(i_clk), .Q(n_0_12), .QN());
   DFF_X1 \b_reg[16]  (.D(i_b[16]), .CK(i_clk), .Q(n_0_13), .QN());
   DFF_X1 \b_reg[15]  (.D(i_b[15]), .CK(i_clk), .Q(n_0_14), .QN());
   DFF_X1 \b_reg[14]  (.D(i_b[14]), .CK(i_clk), .Q(n_0_15), .QN());
   DFF_X1 \b_reg[13]  (.D(i_b[13]), .CK(i_clk), .Q(n_0_16), .QN());
   DFF_X1 \b_reg[12]  (.D(i_b[12]), .CK(i_clk), .Q(n_0_17), .QN());
   DFF_X1 \b_reg[11]  (.D(i_b[11]), .CK(i_clk), .Q(n_0_18), .QN());
   DFF_X1 \b_reg[10]  (.D(i_b[10]), .CK(i_clk), .Q(n_0_19), .QN());
   DFF_X1 \b_reg[9]  (.D(i_b[9]), .CK(i_clk), .Q(n_0_20), .QN());
   DFF_X1 \b_reg[8]  (.D(i_b[8]), .CK(i_clk), .Q(n_0_21), .QN());
   DFF_X1 \b_reg[7]  (.D(i_b[7]), .CK(i_clk), .Q(n_0_22), .QN());
   DFF_X1 \b_reg[6]  (.D(i_b[6]), .CK(i_clk), .Q(n_0_23), .QN());
   DFF_X1 \b_reg[5]  (.D(i_b[5]), .CK(i_clk), .Q(n_0_24), .QN());
   DFF_X1 \b_reg[4]  (.D(i_b[4]), .CK(i_clk), .Q(n_0_25), .QN());
   DFF_X1 \b_reg[3]  (.D(i_b[3]), .CK(i_clk), .Q(n_0_26), .QN());
   DFF_X1 \b_reg[2]  (.D(i_b[2]), .CK(i_clk), .Q(n_0_27), .QN());
   DFF_X1 \b_reg[1]  (.D(i_b[1]), .CK(i_clk), .Q(n_0_28), .QN());
   DFF_X1 \b_reg[0]  (.D(i_b[0]), .CK(i_clk), .Q(n_0_29), .QN());
   DFF_X1 \a_reg[31]  (.D(i_a[31]), .CK(i_clk), .Q(Sa), .QN());
   DFF_X1 \a_reg[30]  (.D(i_a[30]), .CK(i_clk), .Q(n_0_30), .QN());
   DFF_X1 \a_reg[29]  (.D(i_a[29]), .CK(i_clk), .Q(n_0_31), .QN());
   DFF_X1 \a_reg[28]  (.D(i_a[28]), .CK(i_clk), .Q(n_0_32), .QN());
   DFF_X1 \a_reg[27]  (.D(i_a[27]), .CK(i_clk), .Q(n_0_33), .QN());
   DFF_X1 \a_reg[26]  (.D(i_a[26]), .CK(i_clk), .Q(n_0_34), .QN());
   DFF_X1 \a_reg[25]  (.D(i_a[25]), .CK(i_clk), .Q(n_0_35), .QN());
   DFF_X1 \a_reg[24]  (.D(i_a[24]), .CK(i_clk), .Q(n_0_36), .QN());
   DFF_X1 \a_reg[23]  (.D(i_a[23]), .CK(i_clk), .Q(n_0_37), .QN());
   DFF_X1 \a_reg[22]  (.D(i_a[22]), .CK(i_clk), .Q(n_0_38), .QN());
   DFF_X1 \a_reg[21]  (.D(i_a[21]), .CK(i_clk), .Q(n_0_39), .QN());
   DFF_X1 \a_reg[20]  (.D(i_a[20]), .CK(i_clk), .Q(n_0_40), .QN());
   DFF_X1 \a_reg[19]  (.D(i_a[19]), .CK(i_clk), .Q(n_0_41), .QN());
   DFF_X1 \a_reg[18]  (.D(i_a[18]), .CK(i_clk), .Q(n_0_42), .QN());
   DFF_X1 \a_reg[17]  (.D(i_a[17]), .CK(i_clk), .Q(n_0_43), .QN());
   DFF_X1 \a_reg[16]  (.D(i_a[16]), .CK(i_clk), .Q(n_0_44), .QN());
   DFF_X1 \a_reg[15]  (.D(i_a[15]), .CK(i_clk), .Q(n_0_45), .QN());
   DFF_X1 \a_reg[14]  (.D(i_a[14]), .CK(i_clk), .Q(n_0_46), .QN());
   DFF_X1 \a_reg[13]  (.D(i_a[13]), .CK(i_clk), .Q(n_0_47), .QN());
   DFF_X1 \a_reg[12]  (.D(i_a[12]), .CK(i_clk), .Q(n_0_48), .QN());
   DFF_X1 \a_reg[11]  (.D(i_a[11]), .CK(i_clk), .Q(n_0_49), .QN());
   DFF_X1 \a_reg[10]  (.D(i_a[10]), .CK(i_clk), .Q(n_0_50), .QN());
   DFF_X1 \a_reg[9]  (.D(i_a[9]), .CK(i_clk), .Q(n_0_51), .QN());
   DFF_X1 \a_reg[8]  (.D(i_a[8]), .CK(i_clk), .Q(n_0_52), .QN());
   DFF_X1 \a_reg[7]  (.D(i_a[7]), .CK(i_clk), .Q(n_0_53), .QN());
   DFF_X1 \a_reg[6]  (.D(i_a[6]), .CK(i_clk), .Q(n_0_54), .QN());
   DFF_X1 \a_reg[5]  (.D(i_a[5]), .CK(i_clk), .Q(n_0_55), .QN());
   DFF_X1 \a_reg[4]  (.D(i_a[4]), .CK(i_clk), .Q(n_0_56), .QN());
   DFF_X1 \a_reg[3]  (.D(i_a[3]), .CK(i_clk), .Q(n_0_57), .QN());
   DFF_X1 \a_reg[2]  (.D(i_a[2]), .CK(i_clk), .Q(n_0_58), .QN());
   DFF_X1 \a_reg[1]  (.D(i_a[1]), .CK(i_clk), .Q(n_0_59), .QN());
   DFF_X1 \a_reg[0]  (.D(i_a[0]), .CK(i_clk), .Q(n_0_60), .QN());
   FA_X1 i_0_0_0 (.A(mult_res[47]), .B(n_0_0_34), .CI(Eb[0]), .CO(n_0_0_0), 
      .S(E_sum[0]));
   FA_X1 i_0_0_1 (.A(Eb[1]), .B(n_0_0_32), .CI(n_0_0_0), .CO(n_0_0_1), .S(
      E_sum[1]));
   FA_X1 i_0_0_2 (.A(Eb[2]), .B(n_0_0_30), .CI(n_0_0_1), .CO(n_0_0_2), .S(
      E_sum[2]));
   FA_X1 i_0_0_3 (.A(Eb[3]), .B(n_0_0_99), .CI(n_0_0_2), .CO(n_0_0_3), .S(
      E_sum[3]));
   FA_X1 i_0_0_4 (.A(Eb[4]), .B(n_0_0_25), .CI(n_0_0_3), .CO(n_0_0_4), .S(
      E_sum[4]));
   FA_X1 i_0_0_5 (.A(Eb[5]), .B(n_0_0_23), .CI(n_0_0_4), .CO(n_0_0_5), .S(
      E_sum[5]));
   FA_X1 i_0_0_6 (.A(Eb[6]), .B(n_0_0_21), .CI(n_0_0_5), .CO(n_0_0_6), .S(
      E_sum[6]));
   FA_X1 i_0_0_7 (.A(Eb[7]), .B(n_0_0_19), .CI(n_0_0_6), .CO(E_sum[8]), .S(
      E_sum[7]));
   HA_X1 i_0_0_8 (.A(E_sum[1]), .B(E_sum[0]), .CO(n_0_0_7), .S(n_0_0_12));
   HA_X1 i_0_0_9 (.A(E_sum[2]), .B(n_0_0_7), .CO(n_0_0_8), .S(n_0_0_13));
   HA_X1 i_0_0_10 (.A(E_sum[3]), .B(n_0_0_8), .CO(n_0_0_9), .S(n_0_0_14));
   HA_X1 i_0_0_11 (.A(E_sum[4]), .B(n_0_0_9), .CO(n_0_0_10), .S(n_0_0_15));
   HA_X1 i_0_0_12 (.A(E_sum[5]), .B(n_0_0_10), .CO(n_0_0_11), .S(n_0_0_16));
   HA_X1 i_0_0_13 (.A(E_sum[6]), .B(n_0_0_11), .CO(n_0_0_18), .S(n_0_0_17));
   OAI21_X1 i_0_0_14 (.A(n_0_0_113), .B1(n_0_0_119), .B2(n_0_0_118), .ZN(
      n_0_0_19));
   INV_X1 i_0_0_15 (.A(n_0_0_20), .ZN(Eb[7]));
   AOI22_X1 i_0_0_16 (.A1(n_0_0), .A2(n_0_0_73), .B1(n_0_30), .B2(n_0_0_63), 
      .ZN(n_0_0_20));
   OAI21_X1 i_0_0_17 (.A(n_0_0_120), .B1(n_0_0_127), .B2(n_0_0_121), .ZN(
      n_0_0_21));
   INV_X1 i_0_0_18 (.A(n_0_0_22), .ZN(Eb[6]));
   AOI22_X1 i_0_0_19 (.A1(n_0_1), .A2(n_0_0_73), .B1(n_0_31), .B2(n_0_0_63), 
      .ZN(n_0_0_22));
   OAI21_X1 i_0_0_20 (.A(n_0_0_128), .B1(n_0_0_134), .B2(n_0_0_129), .ZN(
      n_0_0_23));
   INV_X1 i_0_0_21 (.A(n_0_0_24), .ZN(Eb[5]));
   AOI22_X1 i_0_0_22 (.A1(n_0_2), .A2(n_0_0_73), .B1(n_0_32), .B2(n_0_0_63), 
      .ZN(n_0_0_24));
   XOR2_X1 i_0_0_23 (.A(n_0_0_147), .B(n_0_0_26), .Z(n_0_0_25));
   AOI21_X1 i_0_0_24 (.A(n_0_0_154), .B1(shamt[4]), .B2(n_0_0_175), .ZN(n_0_0_26));
   INV_X1 i_0_0_25 (.A(n_0_0_27), .ZN(Eb[4]));
   AOI22_X1 i_0_0_26 (.A1(n_0_3), .A2(n_0_0_73), .B1(n_0_33), .B2(n_0_0_63), 
      .ZN(n_0_0_27));
   INV_X1 i_0_0_27 (.A(n_0_0_29), .ZN(Eb[3]));
   AOI22_X1 i_0_0_28 (.A1(n_0_4), .A2(n_0_0_73), .B1(n_0_34), .B2(n_0_0_63), 
      .ZN(n_0_0_29));
   XNOR2_X1 i_0_0_30 (.A(n_0_0_75), .B(n_0_0_89), .ZN(n_0_0_30));
   INV_X1 i_0_0_31 (.A(n_0_0_31), .ZN(Eb[2]));
   AOI22_X1 i_0_0_32 (.A1(n_0_5), .A2(n_0_0_73), .B1(n_0_35), .B2(n_0_0_63), 
      .ZN(n_0_0_31));
   XNOR2_X1 i_0_0_33 (.A(n_0_0_85), .B(n_0_0_88), .ZN(n_0_0_32));
   INV_X1 i_0_0_34 (.A(n_0_0_33), .ZN(Eb[1]));
   AOI22_X1 i_0_0_35 (.A1(n_0_6), .A2(n_0_0_73), .B1(n_0_36), .B2(n_0_0_63), 
      .ZN(n_0_0_33));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_76), .A2(n_0_69), .ZN(Eb[0]));
   OAI21_X1 i_0_0_37 (.A(n_0_0_85), .B1(shamt[0]), .B2(n_0_0_81), .ZN(n_0_0_34));
   INV_X1 i_0_0_39 (.A(n_0_0_35), .ZN(Na[0]));
   AOI22_X1 i_0_0_40 (.A1(n_0_60), .A2(n_0_0_73), .B1(n_0_29), .B2(n_0_0_63), 
      .ZN(n_0_0_35));
   INV_X1 i_0_0_41 (.A(n_0_0_36), .ZN(Na[1]));
   AOI22_X1 i_0_0_42 (.A1(n_0_59), .A2(n_0_0_73), .B1(n_0_28), .B2(n_0_0_63), 
      .ZN(n_0_0_36));
   INV_X1 i_0_0_43 (.A(n_0_0_37), .ZN(Na[2]));
   AOI22_X1 i_0_0_44 (.A1(n_0_58), .A2(n_0_0_73), .B1(n_0_27), .B2(n_0_0_63), 
      .ZN(n_0_0_37));
   INV_X1 i_0_0_45 (.A(n_0_0_38), .ZN(Na[3]));
   AOI22_X1 i_0_0_46 (.A1(n_0_57), .A2(n_0_0_73), .B1(n_0_26), .B2(n_0_0_63), 
      .ZN(n_0_0_38));
   INV_X1 i_0_0_47 (.A(n_0_0_39), .ZN(Na[4]));
   AOI22_X1 i_0_0_48 (.A1(n_0_56), .A2(n_0_0_73), .B1(n_0_25), .B2(n_0_0_63), 
      .ZN(n_0_0_39));
   INV_X1 i_0_0_49 (.A(n_0_0_40), .ZN(Na[5]));
   AOI22_X1 i_0_0_50 (.A1(n_0_55), .A2(n_0_0_73), .B1(n_0_24), .B2(n_0_0_63), 
      .ZN(n_0_0_40));
   INV_X1 i_0_0_51 (.A(n_0_0_41), .ZN(Na[6]));
   AOI22_X1 i_0_0_52 (.A1(n_0_54), .A2(n_0_0_73), .B1(n_0_23), .B2(n_0_0_63), 
      .ZN(n_0_0_41));
   INV_X1 i_0_0_53 (.A(n_0_0_42), .ZN(Na[7]));
   AOI22_X1 i_0_0_54 (.A1(n_0_53), .A2(n_0_0_73), .B1(n_0_22), .B2(n_0_0_63), 
      .ZN(n_0_0_42));
   INV_X1 i_0_0_55 (.A(n_0_0_43), .ZN(Na[8]));
   AOI22_X1 i_0_0_56 (.A1(n_0_52), .A2(n_0_0_73), .B1(n_0_21), .B2(n_0_0_63), 
      .ZN(n_0_0_43));
   INV_X1 i_0_0_57 (.A(n_0_0_44), .ZN(Na[9]));
   AOI22_X1 i_0_0_58 (.A1(n_0_51), .A2(n_0_0_73), .B1(n_0_20), .B2(n_0_0_63), 
      .ZN(n_0_0_44));
   INV_X1 i_0_0_59 (.A(n_0_0_45), .ZN(Na[10]));
   AOI22_X1 i_0_0_60 (.A1(n_0_50), .A2(n_0_0_73), .B1(n_0_19), .B2(n_0_0_63), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_61 (.A(n_0_0_46), .ZN(Na[11]));
   AOI22_X1 i_0_0_62 (.A1(n_0_49), .A2(n_0_0_73), .B1(n_0_18), .B2(n_0_0_63), 
      .ZN(n_0_0_46));
   INV_X1 i_0_0_63 (.A(n_0_0_47), .ZN(Na[12]));
   AOI22_X1 i_0_0_64 (.A1(n_0_48), .A2(n_0_0_73), .B1(n_0_17), .B2(n_0_0_63), 
      .ZN(n_0_0_47));
   INV_X1 i_0_0_65 (.A(n_0_0_48), .ZN(Na[13]));
   AOI22_X1 i_0_0_66 (.A1(n_0_47), .A2(n_0_0_73), .B1(n_0_16), .B2(n_0_0_63), 
      .ZN(n_0_0_48));
   INV_X1 i_0_0_67 (.A(n_0_0_49), .ZN(Na[14]));
   AOI22_X1 i_0_0_68 (.A1(n_0_46), .A2(n_0_0_73), .B1(n_0_15), .B2(n_0_0_63), 
      .ZN(n_0_0_49));
   INV_X1 i_0_0_69 (.A(n_0_0_50), .ZN(Na[15]));
   AOI22_X1 i_0_0_70 (.A1(n_0_45), .A2(n_0_0_73), .B1(n_0_14), .B2(n_0_0_63), 
      .ZN(n_0_0_50));
   INV_X1 i_0_0_71 (.A(n_0_0_51), .ZN(Na[16]));
   AOI22_X1 i_0_0_72 (.A1(n_0_44), .A2(n_0_0_73), .B1(n_0_13), .B2(n_0_0_63), 
      .ZN(n_0_0_51));
   INV_X1 i_0_0_73 (.A(n_0_0_52), .ZN(Na[17]));
   AOI22_X1 i_0_0_74 (.A1(n_0_43), .A2(n_0_0_73), .B1(n_0_12), .B2(n_0_0_63), 
      .ZN(n_0_0_52));
   INV_X1 i_0_0_75 (.A(n_0_0_53), .ZN(Na[18]));
   AOI22_X1 i_0_0_76 (.A1(n_0_42), .A2(n_0_0_73), .B1(n_0_11), .B2(n_0_0_63), 
      .ZN(n_0_0_53));
   INV_X1 i_0_0_77 (.A(n_0_0_54), .ZN(Na[19]));
   AOI22_X1 i_0_0_78 (.A1(n_0_41), .A2(n_0_0_73), .B1(n_0_10), .B2(n_0_0_63), 
      .ZN(n_0_0_54));
   INV_X1 i_0_0_79 (.A(n_0_0_55), .ZN(Na[20]));
   AOI22_X1 i_0_0_80 (.A1(n_0_40), .A2(n_0_0_73), .B1(n_0_9), .B2(n_0_0_63), 
      .ZN(n_0_0_55));
   INV_X1 i_0_0_81 (.A(n_0_0_56), .ZN(Na[21]));
   AOI22_X1 i_0_0_82 (.A1(n_0_39), .A2(n_0_0_73), .B1(n_0_8), .B2(n_0_0_63), 
      .ZN(n_0_0_56));
   INV_X1 i_0_0_83 (.A(n_0_0_57), .ZN(Na[22]));
   AOI22_X1 i_0_0_84 (.A1(n_0_38), .A2(n_0_0_73), .B1(n_0_7), .B2(n_0_0_63), 
      .ZN(n_0_0_57));
   NAND2_X1 i_0_0_85 (.A1(n_0_0_63), .A2(n_0_0_78), .ZN(Na[23]));
   NAND3_X1 i_0_0_36 (.A1(n_0_0_59), .A2(n_0_0_58), .A3(n_0_0_286), .ZN(res[0]));
   AOI22_X1 i_0_0_38 (.A1(mult_res[24]), .A2(n_0_0_233), .B1(mult_res[23]), 
      .B2(n_0_0_234), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_86 (.A1(n_0_0_330), .A2(n_0_0_60), .ZN(n_0_0_59));
   AOI21_X1 i_0_0_87 (.A(n_0_0_61), .B1(E_sum[0]), .B2(n_0_0_68), .ZN(n_0_0_60));
   AOI221_X1 i_0_0_88 (.A(E_sum[0]), .B1(n_0_0_273), .B2(n_0_0_62), .C1(
      n_0_0_274), .C2(n_0_0_249), .ZN(n_0_0_61));
   AOI22_X1 i_0_0_89 (.A1(n_0_0_64), .A2(n_0_0_218), .B1(n_0_0_225), .B2(
      n_0_0_271), .ZN(n_0_0_62));
   OAI221_X1 i_0_0_90 (.A(n_0_0_223), .B1(mult_res[23]), .B2(n_0_0_220), 
      .C1(mult_res[39]), .C2(n_0_0_289), .ZN(n_0_0_64));
   NAND2_X1 i_0_0_91 (.A1(n_0_0_66), .A2(n_0_0_65), .ZN(res[1]));
   AOI22_X1 i_0_0_92 (.A1(mult_res[24]), .A2(n_0_0_234), .B1(mult_res[25]), 
      .B2(n_0_0_233), .ZN(n_0_0_65));
   AOI21_X1 i_0_0_93 (.A(n_0_0_370), .B1(n_0_0_330), .B2(n_0_0_67), .ZN(n_0_0_66));
   OAI22_X1 i_0_0_94 (.A1(n_0_0_208), .A2(n_0_0_248), .B1(E_sum[0]), .B2(
      n_0_0_68), .ZN(n_0_0_67));
   AOI21_X1 i_0_0_95 (.A(n_0_0_69), .B1(n_0_0_274), .B2(n_0_0_241), .ZN(n_0_0_68));
   AOI221_X1 i_0_0_96 (.A(n_0_0_274), .B1(n_0_0_225), .B2(n_0_0_238), .C1(
      n_0_0_287), .C2(n_0_0_70), .ZN(n_0_0_69));
   AOI21_X1 i_0_0_97 (.A(n_0_0_71), .B1(mult_res[32]), .B2(n_0_0_219), .ZN(
      n_0_0_70));
   NOR2_X1 i_0_0_98 (.A1(n_0_0_222), .A2(n_0_0_72), .ZN(n_0_0_71));
   AOI22_X1 i_0_0_99 (.A1(mult_res[24]), .A2(n_0_0_289), .B1(mult_res[40]), 
      .B2(n_0_0_220), .ZN(n_0_0_72));
   NAND2_X1 i_0_0_100 (.A1(n_0_0_286), .A2(n_0_0_82), .ZN(res[3]));
   AOI222_X1 i_0_0_101 (.A1(mult_res[26]), .A2(n_0_0_234), .B1(mult_res[27]), 
      .B2(n_0_0_233), .C1(n_0_0_330), .C2(n_0_0_83), .ZN(n_0_0_82));
   OAI22_X1 i_0_0_102 (.A1(n_0_0_208), .A2(n_0_0_92), .B1(E_sum[0]), .B2(
      n_0_0_84), .ZN(n_0_0_83));
   AOI22_X1 i_0_0_103 (.A1(n_0_0_273), .A2(n_0_0_241), .B1(E_sum[1]), .B2(
      n_0_0_237), .ZN(n_0_0_84));
   NAND2_X1 i_0_0_104 (.A1(n_0_0_286), .A2(n_0_0_90), .ZN(res[4]));
   AOI221_X1 i_0_0_105 (.A(n_0_0_91), .B1(mult_res[27]), .B2(n_0_0_234), 
      .C1(mult_res[28]), .C2(n_0_0_233), .ZN(n_0_0_90));
   AOI221_X1 i_0_0_106 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_326), .C1(
      n_0_0_208), .C2(n_0_0_92), .ZN(n_0_0_91));
   OAI21_X1 i_0_0_107 (.A(n_0_0_93), .B1(n_0_0_273), .B2(n_0_0_305), .ZN(
      n_0_0_92));
   NAND2_X1 i_0_0_108 (.A1(n_0_0_273), .A2(n_0_0_256), .ZN(n_0_0_93));
   NAND3_X1 i_0_0_109 (.A1(n_0_0_286), .A2(n_0_0_106), .A3(n_0_0_105), .ZN(
      res[6]));
   AOI22_X1 i_0_0_110 (.A1(mult_res[30]), .A2(n_0_0_233), .B1(mult_res[29]), 
      .B2(n_0_0_234), .ZN(n_0_0_105));
   NAND2_X1 i_0_0_111 (.A1(n_0_0_330), .A2(n_0_0_107), .ZN(n_0_0_106));
   AOI22_X1 i_0_0_112 (.A1(E_sum[0]), .A2(n_0_0_117), .B1(n_0_0_208), .B2(
      n_0_0_298), .ZN(n_0_0_107));
   NAND2_X1 i_0_0_113 (.A1(n_0_0_115), .A2(n_0_0_114), .ZN(res[7]));
   AOI21_X1 i_0_0_114 (.A(n_0_0_370), .B1(mult_res[31]), .B2(n_0_0_233), 
      .ZN(n_0_0_114));
   AOI21_X1 i_0_0_115 (.A(n_0_0_116), .B1(mult_res[30]), .B2(n_0_0_234), 
      .ZN(n_0_0_115));
   AOI221_X1 i_0_0_116 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_125), .C1(
      n_0_0_208), .C2(n_0_0_117), .ZN(n_0_0_116));
   AOI22_X1 i_0_0_117 (.A1(n_0_0_274), .A2(n_0_0_133), .B1(n_0_0_273), .B2(
      n_0_0_327), .ZN(n_0_0_117));
   NAND3_X1 i_0_0_118 (.A1(n_0_0_286), .A2(n_0_0_123), .A3(n_0_0_122), .ZN(
      res[8]));
   AOI22_X1 i_0_0_119 (.A1(mult_res[32]), .A2(n_0_0_233), .B1(mult_res[31]), 
      .B2(n_0_0_234), .ZN(n_0_0_122));
   NAND2_X1 i_0_0_120 (.A1(n_0_0_330), .A2(n_0_0_124), .ZN(n_0_0_123));
   AOI22_X1 i_0_0_121 (.A1(E_sum[0]), .A2(n_0_0_132), .B1(n_0_0_208), .B2(
      n_0_0_125), .ZN(n_0_0_124));
   AOI21_X1 i_0_0_122 (.A(n_0_0_126), .B1(n_0_0_274), .B2(n_0_0_139), .ZN(
      n_0_0_125));
   NOR2_X1 i_0_0_123 (.A1(n_0_0_274), .A2(n_0_0_323), .ZN(n_0_0_126));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_286), .A2(n_0_0_130), .ZN(res[9]));
   AOI221_X1 i_0_0_125 (.A(n_0_0_131), .B1(mult_res[32]), .B2(n_0_0_234), 
      .C1(mult_res[33]), .C2(n_0_0_233), .ZN(n_0_0_130));
   AOI221_X1 i_0_0_126 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_137), .C1(
      n_0_0_208), .C2(n_0_0_132), .ZN(n_0_0_131));
   AOI22_X1 i_0_0_127 (.A1(n_0_0_273), .A2(n_0_0_133), .B1(n_0_0_274), .B2(
      n_0_0_146), .ZN(n_0_0_132));
   OAI22_X1 i_0_0_128 (.A1(n_0_0_225), .A2(n_0_0_240), .B1(n_0_0_287), .B2(
      n_0_0_161), .ZN(n_0_0_133));
   NAND2_X1 i_0_0_129 (.A1(n_0_0_286), .A2(n_0_0_135), .ZN(res[10]));
   AOI221_X1 i_0_0_130 (.A(n_0_0_136), .B1(mult_res[34]), .B2(n_0_0_233), 
      .C1(mult_res[33]), .C2(n_0_0_234), .ZN(n_0_0_135));
   AOI221_X1 i_0_0_131 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_144), .C1(
      n_0_0_208), .C2(n_0_0_137), .ZN(n_0_0_136));
   OAI21_X1 i_0_0_132 (.A(n_0_0_138), .B1(n_0_0_274), .B2(n_0_0_139), .ZN(
      n_0_0_137));
   NAND2_X1 i_0_0_133 (.A1(n_0_0_274), .A2(n_0_0_152), .ZN(n_0_0_138));
   AOI22_X1 i_0_0_134 (.A1(n_0_0_287), .A2(n_0_0_322), .B1(n_0_0_225), .B2(
      n_0_0_169), .ZN(n_0_0_139));
   NAND3_X1 i_0_0_135 (.A1(n_0_0_286), .A2(n_0_0_142), .A3(n_0_0_141), .ZN(
      res[11]));
   AOI22_X1 i_0_0_136 (.A1(mult_res[35]), .A2(n_0_0_233), .B1(mult_res[34]), 
      .B2(n_0_0_234), .ZN(n_0_0_141));
   OAI211_X1 i_0_0_137 (.A(n_0_0_143), .B(n_0_0_330), .C1(n_0_0_208), .C2(
      n_0_0_151), .ZN(n_0_0_142));
   NAND2_X1 i_0_0_138 (.A1(n_0_0_208), .A2(n_0_0_144), .ZN(n_0_0_143));
   OAI21_X1 i_0_0_139 (.A(n_0_0_145), .B1(n_0_0_274), .B2(n_0_0_146), .ZN(
      n_0_0_144));
   NAND2_X1 i_0_0_140 (.A1(n_0_0_274), .A2(n_0_0_159), .ZN(n_0_0_145));
   AOI22_X1 i_0_0_141 (.A1(n_0_0_287), .A2(n_0_0_328), .B1(n_0_0_225), .B2(
      n_0_0_174), .ZN(n_0_0_146));
   NAND3_X1 i_0_0_142 (.A1(n_0_0_286), .A2(n_0_0_149), .A3(n_0_0_148), .ZN(
      res[12]));
   AOI22_X1 i_0_0_143 (.A1(mult_res[36]), .A2(n_0_0_233), .B1(mult_res[35]), 
      .B2(n_0_0_234), .ZN(n_0_0_148));
   OAI21_X1 i_0_0_144 (.A(n_0_0_150), .B1(E_sum[0]), .B2(n_0_0_151), .ZN(
      n_0_0_149));
   AOI21_X1 i_0_0_145 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_157), .ZN(
      n_0_0_150));
   AOI22_X1 i_0_0_146 (.A1(n_0_0_274), .A2(n_0_0_167), .B1(n_0_0_273), .B2(
      n_0_0_152), .ZN(n_0_0_151));
   AOI22_X1 i_0_0_147 (.A1(mult_res[39]), .A2(n_0_0_201), .B1(n_0_0_287), 
      .B2(n_0_0_324), .ZN(n_0_0_152));
   NAND2_X1 i_0_0_148 (.A1(n_0_0_286), .A2(n_0_0_155), .ZN(res[13]));
   AOI221_X1 i_0_0_149 (.A(n_0_0_156), .B1(mult_res[36]), .B2(n_0_0_234), 
      .C1(mult_res[37]), .C2(n_0_0_233), .ZN(n_0_0_155));
   AOI221_X1 i_0_0_150 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_165), .C1(
      n_0_0_208), .C2(n_0_0_157), .ZN(n_0_0_156));
   AOI21_X1 i_0_0_151 (.A(n_0_0_158), .B1(n_0_0_274), .B2(n_0_0_173), .ZN(
      n_0_0_157));
   NOR2_X1 i_0_0_152 (.A1(n_0_0_274), .A2(n_0_0_159), .ZN(n_0_0_158));
   AOI22_X1 i_0_0_153 (.A1(n_0_0_287), .A2(n_0_0_160), .B1(mult_res[40]), 
      .B2(n_0_0_201), .ZN(n_0_0_159));
   INV_X1 i_0_0_154 (.A(n_0_0_161), .ZN(n_0_0_160));
   AOI22_X1 i_0_0_155 (.A1(mult_res[36]), .A2(n_0_0_270), .B1(mult_res[44]), 
      .B2(n_0_0_219), .ZN(n_0_0_161));
   NAND2_X1 i_0_0_156 (.A1(n_0_0_163), .A2(n_0_0_162), .ZN(res[14]));
   AOI21_X1 i_0_0_157 (.A(n_0_0_370), .B1(mult_res[38]), .B2(n_0_0_233), 
      .ZN(n_0_0_162));
   AOI21_X1 i_0_0_158 (.A(n_0_0_164), .B1(mult_res[37]), .B2(n_0_0_234), 
      .ZN(n_0_0_163));
   AOI221_X1 i_0_0_159 (.A(n_0_0_276), .B1(n_0_0_208), .B2(n_0_0_165), .C1(
      E_sum[0]), .C2(n_0_0_172), .ZN(n_0_0_164));
   INV_X1 i_0_0_160 (.A(n_0_0_166), .ZN(n_0_0_165));
   AOI22_X1 i_0_0_161 (.A1(n_0_0_273), .A2(n_0_0_167), .B1(n_0_0_274), .B2(
      n_0_0_182), .ZN(n_0_0_166));
   AOI22_X1 i_0_0_162 (.A1(n_0_0_287), .A2(n_0_0_168), .B1(mult_res[41]), 
      .B2(n_0_0_201), .ZN(n_0_0_167));
   INV_X1 i_0_0_163 (.A(n_0_0_169), .ZN(n_0_0_168));
   AOI22_X1 i_0_0_164 (.A1(mult_res[37]), .A2(n_0_0_270), .B1(mult_res[45]), 
      .B2(n_0_0_219), .ZN(n_0_0_169));
   NAND2_X1 i_0_0_165 (.A1(n_0_0_286), .A2(n_0_0_170), .ZN(res[15]));
   AOI221_X1 i_0_0_166 (.A(n_0_0_171), .B1(mult_res[38]), .B2(n_0_0_234), 
      .C1(mult_res[39]), .C2(n_0_0_233), .ZN(n_0_0_170));
   AOI221_X1 i_0_0_167 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_180), .C1(
      n_0_0_208), .C2(n_0_0_172), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_168 (.A1(n_0_0_274), .A2(n_0_0_188), .B1(n_0_0_273), .B2(
      n_0_0_173), .ZN(n_0_0_172));
   OAI21_X1 i_0_0_169 (.A(n_0_0_176), .B1(n_0_0_225), .B2(n_0_0_174), .ZN(
      n_0_0_173));
   AOI22_X1 i_0_0_170 (.A1(mult_res[38]), .A2(n_0_0_270), .B1(mult_res[46]), 
      .B2(n_0_0_219), .ZN(n_0_0_174));
   NAND2_X1 i_0_0_171 (.A1(mult_res[42]), .A2(n_0_0_201), .ZN(n_0_0_176));
   NAND2_X1 i_0_0_221 (.A1(n_0_0_178), .A2(n_0_0_177), .ZN(res[16]));
   AOI21_X1 i_0_0_222 (.A(n_0_0_370), .B1(mult_res[40]), .B2(n_0_0_233), 
      .ZN(n_0_0_177));
   AOI21_X1 i_0_0_223 (.A(n_0_0_179), .B1(mult_res[39]), .B2(n_0_0_234), 
      .ZN(n_0_0_178));
   AOI221_X1 i_0_0_224 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_186), .C1(
      n_0_0_208), .C2(n_0_0_180), .ZN(n_0_0_179));
   INV_X1 i_0_0_172 (.A(n_0_0_181), .ZN(n_0_0_180));
   AOI22_X1 i_0_0_173 (.A1(n_0_0_273), .A2(n_0_0_182), .B1(n_0_0_274), .B2(
      n_0_0_195), .ZN(n_0_0_181));
   AOI22_X1 i_0_0_174 (.A1(mult_res[39]), .A2(n_0_0_341), .B1(mult_res[43]), 
      .B2(n_0_0_201), .ZN(n_0_0_182));
   NAND2_X1 i_0_0_228 (.A1(n_0_0_184), .A2(n_0_0_183), .ZN(res[17]));
   AOI21_X1 i_0_0_229 (.A(n_0_0_370), .B1(mult_res[41]), .B2(n_0_0_233), 
      .ZN(n_0_0_183));
   AOI21_X1 i_0_0_230 (.A(n_0_0_185), .B1(mult_res[40]), .B2(n_0_0_234), 
      .ZN(n_0_0_184));
   AOI221_X1 i_0_0_231 (.A(n_0_0_276), .B1(n_0_0_208), .B2(n_0_0_186), .C1(
      E_sum[0]), .C2(n_0_0_192), .ZN(n_0_0_185));
   OAI21_X1 i_0_0_232 (.A(n_0_0_187), .B1(n_0_0_274), .B2(n_0_0_188), .ZN(
      n_0_0_186));
   NAND2_X1 i_0_0_233 (.A1(n_0_0_274), .A2(n_0_0_200), .ZN(n_0_0_187));
   INV_X1 i_0_0_175 (.A(n_0_0_189), .ZN(n_0_0_188));
   AOI22_X1 i_0_0_176 (.A1(mult_res[40]), .A2(n_0_0_341), .B1(mult_res[44]), 
      .B2(n_0_0_201), .ZN(n_0_0_189));
   NAND3_X1 i_0_0_236 (.A1(n_0_0_286), .A2(n_0_0_191), .A3(n_0_0_190), .ZN(
      res[18]));
   AOI22_X1 i_0_0_237 (.A1(mult_res[42]), .A2(n_0_0_233), .B1(mult_res[41]), 
      .B2(n_0_0_234), .ZN(n_0_0_190));
   OAI221_X1 i_0_0_238 (.A(n_0_0_330), .B1(E_sum[0]), .B2(n_0_0_193), .C1(
      n_0_0_208), .C2(n_0_0_198), .ZN(n_0_0_191));
   INV_X1 i_0_0_239 (.A(n_0_0_193), .ZN(n_0_0_192));
   OAI21_X1 i_0_0_240 (.A(n_0_0_194), .B1(n_0_0_274), .B2(n_0_0_195), .ZN(
      n_0_0_193));
   NAND3_X1 i_0_0_241 (.A1(mult_res[43]), .A2(n_0_0_341), .A3(n_0_0_274), 
      .ZN(n_0_0_194));
   AOI22_X1 i_0_0_177 (.A1(mult_res[41]), .A2(n_0_0_341), .B1(mult_res[45]), 
      .B2(n_0_0_201), .ZN(n_0_0_195));
   OAI211_X1 i_0_0_243 (.A(n_0_0_286), .B(n_0_0_196), .C1(n_0_0_276), .C2(
      n_0_0_197), .ZN(res[19]));
   AOI22_X1 i_0_0_244 (.A1(mult_res[43]), .A2(n_0_0_233), .B1(mult_res[42]), 
      .B2(n_0_0_234), .ZN(n_0_0_196));
   AOI21_X1 i_0_0_245 (.A(n_0_0_202), .B1(n_0_0_208), .B2(n_0_0_198), .ZN(
      n_0_0_197));
   OAI21_X1 i_0_0_246 (.A(n_0_0_199), .B1(n_0_0_274), .B2(n_0_0_200), .ZN(
      n_0_0_198));
   NAND3_X1 i_0_0_247 (.A1(mult_res[44]), .A2(n_0_0_341), .A3(n_0_0_274), 
      .ZN(n_0_0_199));
   AOI22_X1 i_0_0_248 (.A1(mult_res[42]), .A2(n_0_0_341), .B1(mult_res[46]), 
      .B2(n_0_0_201), .ZN(n_0_0_200));
   AND2_X1 i_0_0_178 (.A1(n_0_0_270), .A2(n_0_0_225), .ZN(n_0_0_201));
   AND3_X1 i_0_0_250 (.A1(E_sum[0]), .A2(n_0_0_206), .A3(n_0_0_341), .ZN(
      n_0_0_202));
   NAND2_X1 i_0_0_251 (.A1(n_0_0_210), .A2(n_0_0_203), .ZN(res[20]));
   AOI22_X1 i_0_0_252 (.A1(n_0_0_334), .A2(n_0_0_204), .B1(mult_res[43]), 
      .B2(n_0_0_234), .ZN(n_0_0_203));
   OAI21_X1 i_0_0_253 (.A(n_0_0_205), .B1(n_0_0_208), .B2(n_0_0_209), .ZN(
      n_0_0_204));
   NAND2_X1 i_0_0_254 (.A1(n_0_0_208), .A2(n_0_0_206), .ZN(n_0_0_205));
   AOI22_X1 i_0_0_179 (.A1(n_0_0_292), .A2(n_0_0_273), .B1(n_0_0_347), .B2(
      n_0_0_274), .ZN(n_0_0_206));
   AOI22_X1 i_0_0_258 (.A1(mult_res[46]), .A2(n_0_0_228), .B1(mult_res[44]), 
      .B2(E_sum[1]), .ZN(n_0_0_209));
   AOI21_X1 i_0_0_259 (.A(n_0_0_370), .B1(mult_res[44]), .B2(n_0_0_233), 
      .ZN(n_0_0_210));
   NAND2_X1 i_0_0_180 (.A1(n_0_0_215), .A2(n_0_0_211), .ZN(res[21]));
   AOI22_X1 i_0_0_181 (.A1(mult_res[44]), .A2(n_0_0_234), .B1(n_0_0_334), 
      .B2(n_0_0_212), .ZN(n_0_0_211));
   OAI211_X1 i_0_0_182 (.A(n_0_0_213), .B(n_0_0_214), .C1(n_0_0_293), .C2(
      n_0_0_227), .ZN(n_0_0_212));
   NAND3_X1 i_0_0_183 (.A1(n_0_0_208), .A2(E_sum[1]), .A3(mult_res[46]), 
      .ZN(n_0_0_213));
   NAND2_X1 i_0_0_184 (.A1(mult_res[45]), .A2(n_0_0_275), .ZN(n_0_0_214));
   AOI21_X1 i_0_0_185 (.A(n_0_0_370), .B1(mult_res[45]), .B2(n_0_0_233), 
      .ZN(n_0_0_215));
   NOR2_X1 i_0_0_186 (.A1(n_0_0_295), .A2(n_0_0_111), .ZN(n_0_62));
   INV_X1 i_0_0_187 (.A(n_0_0_257), .ZN(res[23]));
   AOI21_X1 i_0_0_188 (.A(n_0_0_266), .B1(n_0_0_208), .B2(n_0_0_110), .ZN(
      n_0_0_257));
   INV_X1 i_0_0_311 (.A(n_0_0_258), .ZN(res[24]));
   AOI21_X1 i_0_0_312 (.A(n_0_0_266), .B1(n_0_0_12), .B2(n_0_0_110), .ZN(
      n_0_0_258));
   INV_X1 i_0_0_313 (.A(n_0_0_259), .ZN(res[25]));
   AOI21_X1 i_0_0_314 (.A(n_0_0_266), .B1(n_0_0_13), .B2(n_0_0_110), .ZN(
      n_0_0_259));
   INV_X1 i_0_0_315 (.A(n_0_0_260), .ZN(res[26]));
   AOI21_X1 i_0_0_316 (.A(n_0_0_266), .B1(n_0_0_14), .B2(n_0_0_110), .ZN(
      n_0_0_260));
   INV_X1 i_0_0_317 (.A(n_0_0_261), .ZN(res[27]));
   AOI21_X1 i_0_0_318 (.A(n_0_0_266), .B1(n_0_0_15), .B2(n_0_0_110), .ZN(
      n_0_0_261));
   INV_X1 i_0_0_319 (.A(n_0_0_262), .ZN(res[28]));
   AOI21_X1 i_0_0_320 (.A(n_0_0_266), .B1(n_0_0_16), .B2(n_0_0_110), .ZN(
      n_0_0_262));
   INV_X1 i_0_0_321 (.A(n_0_0_263), .ZN(res[29]));
   AOI21_X1 i_0_0_322 (.A(n_0_0_266), .B1(n_0_0_17), .B2(n_0_0_110), .ZN(
      n_0_0_263));
   INV_X1 i_0_0_189 (.A(n_0_0_264), .ZN(res[30]));
   AOI21_X1 i_0_0_190 (.A(n_0_0_266), .B1(n_0_0_110), .B2(n_0_0_104), .ZN(
      n_0_0_264));
   INV_X1 i_0_0_191 (.A(n_0_0_267), .ZN(n_0_0_266));
   AOI22_X1 i_0_0_192 (.A1(special_res[23]), .A2(n_0_0_295), .B1(n_0_0_108), 
      .B2(n_0_0_110), .ZN(n_0_0_267));
   NOR3_X1 i_0_0_193 (.A1(shamt[0]), .A2(n_0_0_382), .A3(n_0_0_380), .ZN(Nb[0]));
   OAI22_X1 i_0_0_194 (.A1(shamt[0]), .A2(n_0_0_301), .B1(n_0_0_377), .B2(
      n_0_0_300), .ZN(Nb[2]));
   NAND2_X1 i_0_0_195 (.A1(shamt[0]), .A2(n_0_0_304), .ZN(n_0_0_300));
   AOI22_X1 i_0_0_196 (.A1(n_0_0_390), .A2(n_0_0_303), .B1(shamt[0]), .B2(
      n_0_0_301), .ZN(Nb[3]));
   AOI22_X1 i_0_0_197 (.A1(n_0_70), .A2(n_0_0_310), .B1(n_0_72), .B2(n_0_0_304), 
      .ZN(n_0_0_301));
   OAI21_X1 i_0_0_198 (.A(n_0_0_302), .B1(n_0_0_390), .B2(n_0_0_303), .ZN(Nb[4]));
   NAND2_X1 i_0_0_199 (.A1(n_0_0_390), .A2(n_0_0_307), .ZN(n_0_0_302));
   AOI22_X1 i_0_0_200 (.A1(n_0_71), .A2(n_0_0_310), .B1(n_0_73), .B2(n_0_0_304), 
      .ZN(n_0_0_303));
   INV_X1 i_0_0_201 (.A(n_0_0_382), .ZN(n_0_0_304));
   INV_X1 i_0_0_202 (.A(n_0_0_306), .ZN(Nb[5]));
   AOI22_X1 i_0_0_203 (.A1(shamt[0]), .A2(n_0_0_307), .B1(n_0_0_390), .B2(
      n_0_0_309), .ZN(n_0_0_306));
   OAI22_X1 i_0_0_204 (.A1(shamt[1]), .A2(n_0_0_314), .B1(n_0_0_415), .B2(
      n_0_0_311), .ZN(n_0_0_307));
   INV_X1 i_0_0_205 (.A(n_0_0_308), .ZN(Nb[6]));
   AOI22_X1 i_0_0_206 (.A1(shamt[0]), .A2(n_0_0_309), .B1(n_0_0_390), .B2(
      n_0_0_313), .ZN(n_0_0_308));
   OAI22_X1 i_0_0_207 (.A1(shamt[1]), .A2(n_0_0_317), .B1(n_0_0_416), .B2(
      n_0_0_311), .ZN(n_0_0_309));
   INV_X1 i_0_0_208 (.A(n_0_0_311), .ZN(n_0_0_310));
   NAND2_X1 i_0_0_209 (.A1(shamt[1]), .A2(n_0_0_386), .ZN(n_0_0_311));
   INV_X1 i_0_0_210 (.A(n_0_0_312), .ZN(Nb[7]));
   AOI22_X1 i_0_0_211 (.A1(shamt[0]), .A2(n_0_0_313), .B1(n_0_0_390), .B2(
      n_0_0_316), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_212 (.A1(n_0_0_393), .A2(n_0_0_314), .B1(shamt[1]), .B2(
      n_0_0_321), .ZN(n_0_0_313));
   AOI22_X1 i_0_0_213 (.A1(n_0_70), .A2(n_0_0_424), .B1(n_0_74), .B2(n_0_0_386), 
      .ZN(n_0_0_314));
   INV_X1 i_0_0_214 (.A(n_0_0_315), .ZN(Nb[8]));
   AOI22_X1 i_0_0_215 (.A1(shamt[0]), .A2(n_0_0_316), .B1(n_0_0_390), .B2(
      n_0_0_319), .ZN(n_0_0_315));
   OAI22_X1 i_0_0_216 (.A1(n_0_0_393), .A2(n_0_0_317), .B1(shamt[1]), .B2(
      n_0_0_410), .ZN(n_0_0_316));
   AOI22_X1 i_0_0_217 (.A1(n_0_71), .A2(n_0_0_424), .B1(n_0_0_386), .B2(n_0_75), 
      .ZN(n_0_0_317));
   INV_X1 i_0_0_218 (.A(n_0_0_318), .ZN(Nb[9]));
   AOI22_X1 i_0_0_219 (.A1(shamt[0]), .A2(n_0_0_319), .B1(n_0_0_390), .B2(
      n_0_0_409), .ZN(n_0_0_318));
   OAI21_X1 i_0_0_220 (.A(n_0_0_320), .B1(n_0_0_393), .B2(n_0_0_321), .ZN(
      n_0_0_319));
   NAND2_X1 i_0_0_225 (.A1(n_0_0_393), .A2(n_0_0_404), .ZN(n_0_0_320));
   AOI22_X1 i_0_0_226 (.A1(n_0_72), .A2(n_0_0_424), .B1(n_0_76), .B2(n_0_0_386), 
      .ZN(n_0_0_321));
   OAI22_X1 i_0_0_227 (.A1(n_0_0_390), .A2(n_0_0_398), .B1(shamt[0]), .B2(
      n_0_0_329), .ZN(Nb[11]));
   OAI22_X1 i_0_0_234 (.A1(n_0_0_390), .A2(n_0_0_329), .B1(shamt[0]), .B2(
      n_0_0_332), .ZN(Nb[12]));
   AOI22_X1 i_0_0_235 (.A1(shamt[1]), .A2(n_0_0_412), .B1(n_0_0_393), .B2(
      n_0_0_336), .ZN(n_0_0_329));
   OAI22_X1 i_0_0_242 (.A1(n_0_0_390), .A2(n_0_0_332), .B1(shamt[0]), .B2(
      n_0_0_335), .ZN(Nb[13]));
   AOI22_X1 i_0_0_249 (.A1(n_0_0_393), .A2(n_0_0_340), .B1(shamt[1]), .B2(
      n_0_0_400), .ZN(n_0_0_332));
   OAI22_X1 i_0_0_255 (.A1(n_0_0_390), .A2(n_0_0_335), .B1(shamt[0]), .B2(
      n_0_0_339), .ZN(Nb[14]));
   AOI22_X1 i_0_0_256 (.A1(n_0_0_393), .A2(n_0_0_343), .B1(shamt[1]), .B2(
      n_0_0_336), .ZN(n_0_0_335));
   OAI21_X1 i_0_0_257 (.A(n_0_0_337), .B1(shamt[2]), .B2(n_0_0_350), .ZN(
      n_0_0_336));
   NAND2_X1 i_0_0_260 (.A1(n_0_77), .A2(n_0_0_424), .ZN(n_0_0_337));
   OAI22_X1 i_0_0_261 (.A1(n_0_0_390), .A2(n_0_0_339), .B1(shamt[0]), .B2(
      n_0_0_342), .ZN(Nb[15]));
   AOI22_X1 i_0_0_262 (.A1(shamt[1]), .A2(n_0_0_340), .B1(n_0_0_393), .B2(
      n_0_0_346), .ZN(n_0_0_339));
   AOI22_X1 i_0_0_263 (.A1(n_0_0_100), .A2(n_0_0_353), .B1(shamt[2]), .B2(
      n_0_0_407), .ZN(n_0_0_340));
   OAI22_X1 i_0_0_264 (.A1(n_0_0_390), .A2(n_0_0_342), .B1(shamt[0]), .B2(
      n_0_0_345), .ZN(Nb[16]));
   AOI22_X1 i_0_0_265 (.A1(n_0_0_393), .A2(n_0_0_349), .B1(shamt[1]), .B2(
      n_0_0_343), .ZN(n_0_0_342));
   AOI22_X1 i_0_0_266 (.A1(n_0_0_100), .A2(n_0_0_356), .B1(shamt[2]), .B2(
      n_0_0_413), .ZN(n_0_0_343));
   OAI22_X1 i_0_0_267 (.A1(n_0_0_390), .A2(n_0_0_345), .B1(shamt[0]), .B2(
      n_0_0_348), .ZN(Nb[17]));
   AOI22_X1 i_0_0_268 (.A1(n_0_0_393), .A2(n_0_0_352), .B1(shamt[1]), .B2(
      n_0_0_346), .ZN(n_0_0_345));
   AOI22_X1 i_0_0_269 (.A1(n_0_0_100), .A2(n_0_0_359), .B1(shamt[2]), .B2(
      n_0_0_402), .ZN(n_0_0_346));
   OAI22_X1 i_0_0_270 (.A1(n_0_0_390), .A2(n_0_0_348), .B1(shamt[0]), .B2(
      n_0_0_351), .ZN(Nb[18]));
   AOI22_X1 i_0_0_271 (.A1(n_0_0_393), .A2(n_0_0_355), .B1(shamt[1]), .B2(
      n_0_0_349), .ZN(n_0_0_348));
   AOI22_X1 i_0_0_272 (.A1(n_0_0_100), .A2(n_0_0_362), .B1(shamt[2]), .B2(
      n_0_0_350), .ZN(n_0_0_349));
   AOI22_X1 i_0_0_273 (.A1(n_0_0_414), .A2(n_0_73), .B1(n_0_0_425), .B2(n_0_81), 
      .ZN(n_0_0_350));
   OAI22_X1 i_0_0_274 (.A1(n_0_0_390), .A2(n_0_0_351), .B1(shamt[0]), .B2(
      n_0_0_354), .ZN(Nb[19]));
   AOI22_X1 i_0_0_275 (.A1(n_0_0_393), .A2(n_0_0_358), .B1(shamt[1]), .B2(
      n_0_0_352), .ZN(n_0_0_351));
   OAI22_X1 i_0_0_276 (.A1(n_0_0_100), .A2(n_0_0_353), .B1(shamt[2]), .B2(
      n_0_0_395), .ZN(n_0_0_352));
   AOI22_X1 i_0_0_277 (.A1(n_0_0_425), .A2(n_0_82), .B1(n_0_0_414), .B2(n_0_74), 
      .ZN(n_0_0_353));
   OAI22_X1 i_0_0_278 (.A1(n_0_0_390), .A2(n_0_0_354), .B1(shamt[0]), .B2(
      n_0_0_357), .ZN(Nb[20]));
   AOI22_X1 i_0_0_279 (.A1(n_0_0_393), .A2(n_0_0_361), .B1(shamt[1]), .B2(
      n_0_0_355), .ZN(n_0_0_354));
   OAI22_X1 i_0_0_280 (.A1(n_0_0_100), .A2(n_0_0_356), .B1(shamt[2]), .B2(
      n_0_0_379), .ZN(n_0_0_355));
   AOI22_X1 i_0_0_281 (.A1(n_0_0_414), .A2(n_0_75), .B1(n_0_0_425), .B2(n_0_83), 
      .ZN(n_0_0_356));
   OAI22_X1 i_0_0_282 (.A1(n_0_0_390), .A2(n_0_0_357), .B1(shamt[0]), .B2(
      n_0_0_360), .ZN(Nb[21]));
   AOI22_X1 i_0_0_283 (.A1(shamt[1]), .A2(n_0_0_358), .B1(n_0_0_393), .B2(
      n_0_0_389), .ZN(n_0_0_357));
   OAI22_X1 i_0_0_284 (.A1(n_0_0_100), .A2(n_0_0_359), .B1(shamt[2]), .B2(
      n_0_0_399), .ZN(n_0_0_358));
   AOI22_X1 i_0_0_285 (.A1(n_0_84), .A2(n_0_0_425), .B1(n_0_0_414), .B2(n_0_76), 
      .ZN(n_0_0_359));
   OAI22_X1 i_0_0_286 (.A1(n_0_0_390), .A2(n_0_0_360), .B1(shamt[0]), .B2(
      n_0_0_387), .ZN(Nb[22]));
   AOI22_X1 i_0_0_287 (.A1(n_0_0_393), .A2(n_0_0_378), .B1(shamt[1]), .B2(
      n_0_0_361), .ZN(n_0_0_360));
   OAI22_X1 i_0_0_288 (.A1(n_0_0_100), .A2(n_0_0_362), .B1(shamt[2]), .B2(
      n_0_0_368), .ZN(n_0_0_361));
   AOI22_X1 i_0_0_289 (.A1(n_0_0_425), .A2(n_0_85), .B1(n_0_0_414), .B2(n_0_77), 
      .ZN(n_0_0_362));
   OAI21_X1 i_0_0_290 (.A(n_0_0_363), .B1(n_0_0_390), .B2(n_0_0_387), .ZN(Nb[23]));
   OAI21_X1 i_0_0_291 (.A(n_0_0_364), .B1(n_0_0_393), .B2(n_0_0_378), .ZN(
      n_0_0_363));
   AOI21_X1 i_0_0_292 (.A(shamt[0]), .B1(n_0_0_393), .B2(n_0_0_365), .ZN(
      n_0_0_364));
   AOI22_X1 i_0_0_293 (.A1(n_0_0_376), .A2(n_0_0_366), .B1(shamt[2]), .B2(
      n_0_0_367), .ZN(n_0_0_365));
   AOI221_X1 i_0_0_294 (.A(shamt[2]), .B1(n_0_0_425), .B2(n_0_0_372), .C1(
      n_0_0_414), .C2(n_0_0_375), .ZN(n_0_0_366));
   INV_X1 i_0_0_295 (.A(n_0_0_368), .ZN(n_0_0_367));
   AOI222_X1 i_0_0_296 (.A1(n_0_0_405), .A2(n_0_73), .B1(n_0_0_414), .B2(n_0_81), 
      .C1(n_0_0_425), .C2(n_0_65), .ZN(n_0_0_368));
   INV_X1 i_0_0_297 (.A(n_0_0_369), .ZN(n_0_81));
   AOI22_X1 i_0_0_298 (.A1(n_0_18), .A2(n_0_0_73), .B1(n_0_49), .B2(n_0_0_63), 
      .ZN(n_0_0_369));
   INV_X1 i_0_0_299 (.A(n_0_0_371), .ZN(n_0_65));
   AOI22_X1 i_0_0_300 (.A1(n_0_10), .A2(n_0_0_73), .B1(n_0_41), .B2(n_0_0_63), 
      .ZN(n_0_0_371));
   INV_X1 i_0_0_301 (.A(n_0_0_372), .ZN(n_0_69));
   NAND2_X1 i_0_0_302 (.A1(n_0_0_73), .A2(n_0_0_79), .ZN(n_0_0_372));
   INV_X1 i_0_0_303 (.A(n_0_0_375), .ZN(n_0_85));
   AOI22_X1 i_0_0_304 (.A1(n_0_14), .A2(n_0_0_73), .B1(n_0_45), .B2(n_0_0_63), 
      .ZN(n_0_0_375));
   OAI21_X1 i_0_0_305 (.A(shamt[4]), .B1(shamt[3]), .B2(n_0_0_419), .ZN(
      n_0_0_376));
   AOI22_X1 i_0_0_306 (.A1(shamt[2]), .A2(n_0_0_379), .B1(n_0_0_100), .B2(
      n_0_0_383), .ZN(n_0_0_378));
   AOI222_X1 i_0_0_307 (.A1(n_0_0_425), .A2(n_0_63), .B1(n_0_0_414), .B2(n_0_79), 
      .C1(n_0_0_405), .C2(n_0_71), .ZN(n_0_0_379));
   INV_X1 i_0_0_308 (.A(n_0_0_381), .ZN(n_0_63));
   AOI22_X1 i_0_0_309 (.A1(n_0_12), .A2(n_0_0_73), .B1(n_0_43), .B2(n_0_0_63), 
      .ZN(n_0_0_381));
   AOI222_X1 i_0_0_310 (.A1(n_0_0_414), .A2(n_0_83), .B1(n_0_0_425), .B2(n_0_67), 
      .C1(n_0_0_405), .C2(n_0_75), .ZN(n_0_0_383));
   INV_X1 i_0_0_323 (.A(n_0_0_384), .ZN(n_0_67));
   AOI22_X1 i_0_0_324 (.A1(n_0_8), .A2(n_0_0_73), .B1(n_0_39), .B2(n_0_0_63), 
      .ZN(n_0_0_384));
   INV_X1 i_0_0_325 (.A(n_0_0_385), .ZN(n_0_83));
   OAI22_X1 i_0_0_326 (.A1(n_0_47), .A2(n_0_0_73), .B1(n_0_16), .B2(n_0_0_63), 
      .ZN(n_0_0_385));
   AOI21_X1 i_0_0_327 (.A(n_0_0_388), .B1(shamt[1]), .B2(n_0_0_389), .ZN(
      n_0_0_387));
   AOI221_X1 i_0_0_328 (.A(shamt[1]), .B1(n_0_0_100), .B2(n_0_0_403), .C1(
      shamt[2]), .C2(n_0_0_399), .ZN(n_0_0_388));
   OAI22_X1 i_0_0_329 (.A1(n_0_0_100), .A2(n_0_0_395), .B1(shamt[2]), .B2(
      n_0_0_391), .ZN(n_0_0_389));
   AOI222_X1 i_0_0_330 (.A1(n_0_0_414), .A2(n_0_82), .B1(n_0_0_405), .B2(n_0_74), 
      .C1(n_0_0_425), .C2(n_0_66), .ZN(n_0_0_391));
   INV_X1 i_0_0_331 (.A(n_0_0_392), .ZN(n_0_66));
   AOI22_X1 i_0_0_332 (.A1(n_0_9), .A2(n_0_0_73), .B1(n_0_40), .B2(n_0_0_63), 
      .ZN(n_0_0_392));
   INV_X1 i_0_0_333 (.A(n_0_0_394), .ZN(n_0_82));
   AOI22_X1 i_0_0_334 (.A1(n_0_17), .A2(n_0_0_73), .B1(n_0_48), .B2(n_0_0_63), 
      .ZN(n_0_0_394));
   AOI222_X1 i_0_0_335 (.A1(n_0_0_425), .A2(n_0_86), .B1(n_0_0_414), .B2(n_0_78), 
      .C1(n_0_0_405), .C2(n_0_70), .ZN(n_0_0_395));
   INV_X1 i_0_0_336 (.A(n_0_0_397), .ZN(n_0_86));
   AOI22_X1 i_0_0_337 (.A1(n_0_13), .A2(n_0_0_73), .B1(n_0_44), .B2(n_0_0_63), 
      .ZN(n_0_0_397));
   AOI222_X1 i_0_0_338 (.A1(n_0_0_425), .A2(n_0_64), .B1(n_0_0_414), .B2(n_0_80), 
      .C1(n_0_0_405), .C2(n_0_72), .ZN(n_0_0_399));
   INV_X1 i_0_0_339 (.A(n_0_0_401), .ZN(n_0_64));
   AOI22_X1 i_0_0_340 (.A1(n_0_11), .A2(n_0_0_73), .B1(n_0_42), .B2(n_0_0_63), 
      .ZN(n_0_0_401));
   AOI222_X1 i_0_0_341 (.A1(n_0_0_414), .A2(n_0_84), .B1(n_0_0_405), .B2(n_0_76), 
      .C1(n_0_0_425), .C2(n_0_68), .ZN(n_0_0_403));
   NOR2_X1 i_0_0_342 (.A1(n_0_0_428), .A2(shamt[3]), .ZN(n_0_0_405));
   INV_X1 i_0_0_343 (.A(n_0_0_406), .ZN(n_0_68));
   AOI22_X1 i_0_0_344 (.A1(n_0_7), .A2(n_0_0_73), .B1(n_0_38), .B2(n_0_0_63), 
      .ZN(n_0_0_406));
   INV_X1 i_0_0_345 (.A(n_0_0_408), .ZN(n_0_84));
   AOI22_X1 i_0_0_346 (.A1(n_0_15), .A2(n_0_0_73), .B1(n_0_46), .B2(n_0_0_63), 
      .ZN(n_0_0_408));
   INV_X1 i_0_0_347 (.A(outA[0]), .ZN(n_0_0_28));
   NOR3_X1 i_0_0_348 (.A1(n_0_0_28), .A2(outA[1]), .A3(outA[2]), .ZN(n_0_0_63));
   INV_X1 i_0_0_349 (.A(n_0_0_63), .ZN(n_0_0_73));
   AOI22_X1 i_0_0_350 (.A1(n_0_0_73), .A2(n_0_35), .B1(n_0_0_63), .B2(n_0_5), 
      .ZN(n_0_0_74));
   XOR2_X1 i_0_0_351 (.A(n_0_0_74), .B(shamt[2]), .Z(n_0_0_75));
   INV_X1 i_0_0_352 (.A(b), .ZN(n_0_0_76));
   INV_X1 i_0_0_353 (.A(outB[0]), .ZN(n_0_0_77));
   NOR3_X1 i_0_0_354 (.A1(n_0_0_77), .A2(outB[1]), .A3(outB[2]), .ZN(n_0_0_78));
   INV_X1 i_0_0_355 (.A(n_0_0_78), .ZN(n_0_0_79));
   NAND2_X1 i_0_0_356 (.A1(n_0_0_79), .A2(n_0_0_76), .ZN(n_0_0_80));
   AOI22_X1 i_0_0_357 (.A1(n_0_0_73), .A2(n_0_37), .B1(n_0_0_80), .B2(n_0_0_63), 
      .ZN(n_0_0_81));
   NAND2_X1 i_0_0_358 (.A1(n_0_0_81), .A2(shamt[0]), .ZN(n_0_0_85));
   OAI22_X1 i_0_0_359 (.A1(n_0_0_73), .A2(n_0_6), .B1(n_0_0_63), .B2(n_0_36), 
      .ZN(n_0_0_86));
   NAND2_X1 i_0_0_360 (.A1(n_0_0_86), .A2(shamt[1]), .ZN(n_0_0_87));
   OAI21_X1 i_0_0_361 (.A(n_0_0_87), .B1(n_0_0_86), .B2(shamt[1]), .ZN(n_0_0_88));
   OAI21_X1 i_0_0_362 (.A(n_0_0_87), .B1(n_0_0_88), .B2(n_0_0_85), .ZN(n_0_0_89));
   AOI22_X1 i_0_0_363 (.A1(n_0_0_89), .A2(n_0_0_75), .B1(n_0_0_74), .B2(shamt[2]), 
      .ZN(n_0_0_94));
   OAI22_X1 i_0_0_364 (.A1(n_0_0_73), .A2(n_0_4), .B1(n_0_0_63), .B2(n_0_34), 
      .ZN(n_0_0_95));
   OR2_X1 i_0_0_365 (.A1(n_0_0_95), .A2(shamt[3]), .ZN(n_0_0_96));
   NAND2_X1 i_0_0_366 (.A1(n_0_0_95), .A2(shamt[3]), .ZN(n_0_0_97));
   NAND2_X1 i_0_0_367 (.A1(n_0_0_96), .A2(n_0_0_97), .ZN(n_0_0_98));
   XNOR2_X1 i_0_0_368 (.A(n_0_0_94), .B(n_0_0_98), .ZN(n_0_0_99));
   INV_X1 i_0_0_369 (.A(shamt[2]), .ZN(n_0_0_100));
   AND2_X1 i_0_0_370 (.A1(n_0_0_110), .A2(n_0_0_101), .ZN(n_0_61));
   OAI21_X1 i_0_0_371 (.A(n_0_0_109), .B1(n_0_0_103), .B2(n_0_0_102), .ZN(
      n_0_0_101));
   NAND4_X1 i_0_0_372 (.A1(n_0_0_16), .A2(n_0_0_15), .A3(n_0_0_17), .A4(
      n_0_0_104), .ZN(n_0_0_102));
   NAND4_X1 i_0_0_373 (.A1(n_0_0_208), .A2(n_0_0_12), .A3(n_0_0_13), .A4(
      n_0_0_14), .ZN(n_0_0_103));
   OAI21_X1 i_0_0_374 (.A(n_0_0_112), .B1(n_0_0_216), .B2(n_0_0_207), .ZN(
      n_0_0_104));
   INV_X1 i_0_0_375 (.A(n_0_0_109), .ZN(n_0_0_108));
   NAND2_X1 i_0_0_376 (.A1(E_sum[8]), .A2(n_0_0_112), .ZN(n_0_0_109));
   AND3_X1 i_0_0_377 (.A1(enable), .A2(n_0_0_113), .A3(n_0_0_111), .ZN(n_0_0_110));
   NAND3_X1 i_0_0_378 (.A1(n_0_0_216), .A2(n_0_0_207), .A3(n_0_0_217), .ZN(
      n_0_0_111));
   NAND2_X1 i_0_0_379 (.A1(n_0_0_216), .A2(n_0_0_207), .ZN(n_0_0_112));
   NAND2_X1 i_0_0_380 (.A1(n_0_0_119), .A2(n_0_0_118), .ZN(n_0_0_113));
   AOI22_X1 i_0_0_381 (.A1(n_0_0), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_30), 
      .ZN(n_0_0_118));
   INV_X1 i_0_0_382 (.A(n_0_0_120), .ZN(n_0_0_119));
   NAND2_X1 i_0_0_383 (.A1(n_0_0_127), .A2(n_0_0_121), .ZN(n_0_0_120));
   AOI22_X1 i_0_0_384 (.A1(n_0_1), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_31), 
      .ZN(n_0_0_121));
   INV_X1 i_0_0_385 (.A(n_0_0_128), .ZN(n_0_0_127));
   NAND2_X1 i_0_0_386 (.A1(n_0_0_134), .A2(n_0_0_129), .ZN(n_0_0_128));
   AOI22_X1 i_0_0_387 (.A1(n_0_2), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_32), 
      .ZN(n_0_0_129));
   AOI21_X1 i_0_0_388 (.A(n_0_0_154), .B1(n_0_0_147), .B2(n_0_0_140), .ZN(
      n_0_0_134));
   NAND2_X1 i_0_0_389 (.A1(shamt[4]), .A2(n_0_0_175), .ZN(n_0_0_140));
   NAND2_X1 i_0_0_390 (.A1(n_0_0_96), .A2(n_0_0_153), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_391 (.A1(n_0_0_94), .A2(n_0_0_97), .ZN(n_0_0_153));
   NOR2_X1 i_0_0_392 (.A1(shamt[4]), .A2(n_0_0_175), .ZN(n_0_0_154));
   OAI22_X1 i_0_0_393 (.A1(n_0_33), .A2(n_0_0_63), .B1(n_0_3), .B2(n_0_0_73), 
      .ZN(n_0_0_175));
   INV_X1 i_0_0_394 (.A(n_0_0_18), .ZN(n_0_0_207));
   INV_X1 i_0_0_395 (.A(E_sum[0]), .ZN(n_0_0_208));
   INV_X1 i_0_0_396 (.A(E_sum[7]), .ZN(n_0_0_216));
   INV_X1 i_0_0_397 (.A(E_sum[8]), .ZN(n_0_0_217));
   AOI21_X1 i_0_0_398 (.A(n_0_0_225), .B1(mult_res[31]), .B2(n_0_0_219), 
      .ZN(n_0_0_218));
   NOR2_X1 i_0_0_399 (.A1(n_0_0_223), .A2(n_0_0_220), .ZN(n_0_0_219));
   AOI21_X1 i_0_0_400 (.A(n_0_0_221), .B1(E_sum[4]), .B2(n_0_0_224), .ZN(
      n_0_0_220));
   NOR2_X1 i_0_0_401 (.A1(E_sum[4]), .A2(n_0_0_224), .ZN(n_0_0_221));
   INV_X1 i_0_0_402 (.A(n_0_0_223), .ZN(n_0_0_222));
   OAI21_X1 i_0_0_403 (.A(n_0_0_224), .B1(n_0_0_229), .B2(n_0_0_226), .ZN(
      n_0_0_223));
   NAND2_X1 i_0_0_404 (.A1(n_0_0_229), .A2(n_0_0_226), .ZN(n_0_0_224));
   AOI21_X1 i_0_0_405 (.A(n_0_0_226), .B1(E_sum[2]), .B2(n_0_0_227), .ZN(
      n_0_0_225));
   NOR2_X1 i_0_0_406 (.A1(E_sum[2]), .A2(n_0_0_227), .ZN(n_0_0_226));
   NAND2_X1 i_0_0_407 (.A1(n_0_0_228), .A2(n_0_0_208), .ZN(n_0_0_227));
   INV_X1 i_0_0_408 (.A(E_sum[1]), .ZN(n_0_0_228));
   INV_X1 i_0_0_409 (.A(E_sum[3]), .ZN(n_0_0_229));
   NAND2_X1 i_0_0_410 (.A1(n_0_0_286), .A2(n_0_0_230), .ZN(res[2]));
   AOI221_X1 i_0_0_411 (.A(n_0_0_231), .B1(mult_res[26]), .B2(n_0_0_233), 
      .C1(mult_res[25]), .C2(n_0_0_234), .ZN(n_0_0_230));
   AOI211_X1 i_0_0_412 (.A(n_0_0_232), .B(n_0_0_276), .C1(n_0_0_208), .C2(
      n_0_0_248), .ZN(n_0_0_231));
   AOI221_X1 i_0_0_413 (.A(n_0_0_208), .B1(n_0_0_228), .B2(n_0_0_237), .C1(
      n_0_0_273), .C2(n_0_0_241), .ZN(n_0_0_232));
   AND2_X1 i_0_0_414 (.A1(mult_res[47]), .A2(n_0_0_236), .ZN(n_0_0_233));
   NOR2_X1 i_0_0_415 (.A1(mult_res[47]), .A2(n_0_0_235), .ZN(n_0_0_234));
   INV_X1 i_0_0_416 (.A(n_0_0_236), .ZN(n_0_0_235));
   AOI211_X1 i_0_0_417 (.A(n_0_0_282), .B(n_0_0_280), .C1(n_0_0_119), .C2(
      n_0_0_118), .ZN(n_0_0_236));
   AOI22_X1 i_0_0_418 (.A1(n_0_0_287), .A2(n_0_0_238), .B1(n_0_0_225), .B2(
      n_0_0_240), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_419 (.A1(mult_res[36]), .A2(n_0_0_219), .B1(n_0_0_288), 
      .B2(n_0_0_239), .ZN(n_0_0_238));
   OAI22_X1 i_0_0_420 (.A1(n_0_0_291), .A2(n_0_0_220), .B1(n_0_0_293), .B2(
      n_0_0_289), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_421 (.A1(mult_res[32]), .A2(n_0_0_270), .B1(mult_res[40]), 
      .B2(n_0_0_219), .ZN(n_0_0_240));
   OAI22_X1 i_0_0_422 (.A1(n_0_0_225), .A2(n_0_0_242), .B1(n_0_0_287), .B2(
      n_0_0_245), .ZN(n_0_0_241));
   AOI21_X1 i_0_0_423 (.A(n_0_0_243), .B1(mult_res[34]), .B2(n_0_0_219), 
      .ZN(n_0_0_242));
   INV_X1 i_0_0_424 (.A(n_0_0_244), .ZN(n_0_0_243));
   OAI221_X1 i_0_0_425 (.A(n_0_0_223), .B1(mult_res[42]), .B2(n_0_0_289), 
      .C1(mult_res[26]), .C2(n_0_0_220), .ZN(n_0_0_244));
   AOI22_X1 i_0_0_426 (.A1(mult_res[38]), .A2(n_0_0_219), .B1(n_0_0_288), 
      .B2(n_0_0_246), .ZN(n_0_0_245));
   INV_X1 i_0_0_427 (.A(n_0_0_247), .ZN(n_0_0_246));
   OAI22_X1 i_0_0_428 (.A1(mult_res[30]), .A2(n_0_0_220), .B1(mult_res[46]), 
      .B2(n_0_0_289), .ZN(n_0_0_247));
   AOI22_X1 i_0_0_429 (.A1(n_0_0_273), .A2(n_0_0_249), .B1(n_0_0_274), .B2(
      n_0_0_265), .ZN(n_0_0_248));
   OAI22_X1 i_0_0_430 (.A1(n_0_0_225), .A2(n_0_0_250), .B1(n_0_0_287), .B2(
      n_0_0_253), .ZN(n_0_0_249));
   AOI21_X1 i_0_0_431 (.A(n_0_0_251), .B1(mult_res[33]), .B2(n_0_0_219), 
      .ZN(n_0_0_250));
   INV_X1 i_0_0_432 (.A(n_0_0_252), .ZN(n_0_0_251));
   OAI221_X1 i_0_0_433 (.A(n_0_0_223), .B1(mult_res[41]), .B2(n_0_0_289), 
      .C1(mult_res[25]), .C2(n_0_0_220), .ZN(n_0_0_252));
   AOI22_X1 i_0_0_434 (.A1(mult_res[37]), .A2(n_0_0_219), .B1(n_0_0_288), 
      .B2(n_0_0_254), .ZN(n_0_0_253));
   INV_X1 i_0_0_435 (.A(n_0_0_255), .ZN(n_0_0_254));
   OAI22_X1 i_0_0_436 (.A1(mult_res[29]), .A2(n_0_0_220), .B1(mult_res[45]), 
      .B2(n_0_0_289), .ZN(n_0_0_255));
   INV_X1 i_0_0_437 (.A(n_0_0_265), .ZN(n_0_0_256));
   AOI22_X1 i_0_0_438 (.A1(n_0_0_225), .A2(n_0_0_269), .B1(n_0_0_287), .B2(
      n_0_0_271), .ZN(n_0_0_265));
   INV_X1 i_0_0_439 (.A(n_0_0_269), .ZN(n_0_0_268));
   AOI22_X1 i_0_0_440 (.A1(mult_res[31]), .A2(n_0_0_270), .B1(mult_res[39]), 
      .B2(n_0_0_219), .ZN(n_0_0_269));
   NOR2_X1 i_0_0_441 (.A1(n_0_0_220), .A2(n_0_0_222), .ZN(n_0_0_270));
   AOI22_X1 i_0_0_442 (.A1(mult_res[35]), .A2(n_0_0_219), .B1(n_0_0_288), 
      .B2(n_0_0_272), .ZN(n_0_0_271));
   OAI22_X1 i_0_0_443 (.A1(n_0_0_290), .A2(n_0_0_220), .B1(n_0_0_292), .B2(
      n_0_0_289), .ZN(n_0_0_272));
   INV_X1 i_0_0_444 (.A(n_0_0_274), .ZN(n_0_0_273));
   AOI21_X1 i_0_0_445 (.A(n_0_0_275), .B1(n_0_0_208), .B2(n_0_0_228), .ZN(
      n_0_0_274));
   NOR2_X1 i_0_0_446 (.A1(n_0_0_208), .A2(n_0_0_228), .ZN(n_0_0_275));
   NAND4_X1 i_0_0_447 (.A1(n_0_0_113), .A2(n_0_0_277), .A3(n_0_0_279), .A4(
      n_0_0_282), .ZN(n_0_0_276));
   NOR2_X1 i_0_0_448 (.A1(n_0_0_280), .A2(n_0_0_278), .ZN(n_0_0_277));
   AOI22_X1 i_0_0_449 (.A1(n_0_0_294), .A2(n_0_0_221), .B1(E_sum[5]), .B2(
      n_0_0_216), .ZN(n_0_0_278));
   OAI22_X1 i_0_0_450 (.A1(E_sum[5]), .A2(n_0_0_216), .B1(n_0_0_294), .B2(
      n_0_0_221), .ZN(n_0_0_279));
   INV_X1 i_0_0_451 (.A(n_0_0_281), .ZN(n_0_0_280));
   AOI21_X1 i_0_0_452 (.A(n_0_0_295), .B1(n_0_0_111), .B2(n_0_0_101), .ZN(
      n_0_0_281));
   NAND2_X1 i_0_0_453 (.A1(n_0_0_111), .A2(n_0_0_283), .ZN(n_0_0_282));
   NAND3_X1 i_0_0_454 (.A1(n_0_0_285), .A2(n_0_0_284), .A3(n_0_0_217), .ZN(
      n_0_0_283));
   NOR4_X1 i_0_0_455 (.A1(n_0_0_13), .A2(n_0_0_12), .A3(n_0_0_16), .A4(n_0_0_104), 
      .ZN(n_0_0_284));
   NOR4_X1 i_0_0_456 (.A1(n_0_0_208), .A2(n_0_0_14), .A3(n_0_0_15), .A4(n_0_0_17), 
      .ZN(n_0_0_285));
   NAND2_X1 i_0_0_457 (.A1(n_0_0_295), .A2(special_res[0]), .ZN(n_0_0_286));
   INV_X1 i_0_0_458 (.A(n_0_0_225), .ZN(n_0_0_287));
   INV_X1 i_0_0_459 (.A(n_0_0_222), .ZN(n_0_0_288));
   INV_X1 i_0_0_460 (.A(n_0_0_220), .ZN(n_0_0_289));
   INV_X1 i_0_0_461 (.A(mult_res[27]), .ZN(n_0_0_290));
   INV_X1 i_0_0_462 (.A(mult_res[28]), .ZN(n_0_0_291));
   INV_X1 i_0_0_463 (.A(mult_res[43]), .ZN(n_0_0_292));
   INV_X1 i_0_0_464 (.A(mult_res[44]), .ZN(n_0_0_293));
   INV_X1 i_0_0_465 (.A(E_sum[6]), .ZN(n_0_0_294));
   INV_X1 i_0_0_466 (.A(enable), .ZN(n_0_0_295));
   NAND2_X1 i_0_0_467 (.A1(n_0_0_286), .A2(n_0_0_296), .ZN(res[5]));
   AOI221_X1 i_0_0_468 (.A(n_0_0_297), .B1(mult_res[28]), .B2(n_0_0_234), 
      .C1(mult_res[29]), .C2(n_0_0_233), .ZN(n_0_0_296));
   AOI221_X1 i_0_0_469 (.A(n_0_0_276), .B1(E_sum[0]), .B2(n_0_0_298), .C1(
      n_0_0_208), .C2(n_0_0_326), .ZN(n_0_0_297));
   OAI21_X1 i_0_0_470 (.A(n_0_0_299), .B1(n_0_0_274), .B2(n_0_0_305), .ZN(
      n_0_0_298));
   NAND2_X1 i_0_0_471 (.A1(n_0_0_274), .A2(n_0_0_323), .ZN(n_0_0_299));
   AOI22_X1 i_0_0_472 (.A1(n_0_0_287), .A2(n_0_0_253), .B1(n_0_0_225), .B2(
      n_0_0_322), .ZN(n_0_0_305));
   AOI22_X1 i_0_0_473 (.A1(mult_res[33]), .A2(n_0_0_270), .B1(mult_res[41]), 
      .B2(n_0_0_219), .ZN(n_0_0_322));
   AOI22_X1 i_0_0_474 (.A1(n_0_0_287), .A2(n_0_0_268), .B1(n_0_0_225), .B2(
      n_0_0_324), .ZN(n_0_0_323));
   INV_X1 i_0_0_475 (.A(n_0_0_325), .ZN(n_0_0_324));
   AOI22_X1 i_0_0_476 (.A1(mult_res[35]), .A2(n_0_0_270), .B1(mult_res[43]), 
      .B2(n_0_0_219), .ZN(n_0_0_325));
   OAI22_X1 i_0_0_477 (.A1(n_0_0_273), .A2(n_0_0_327), .B1(n_0_0_274), .B2(
      n_0_0_237), .ZN(n_0_0_326));
   OAI22_X1 i_0_0_478 (.A1(n_0_0_287), .A2(n_0_0_328), .B1(n_0_0_225), .B2(
      n_0_0_245), .ZN(n_0_0_327));
   AOI22_X1 i_0_0_479 (.A1(mult_res[34]), .A2(n_0_0_270), .B1(mult_res[42]), 
      .B2(n_0_0_219), .ZN(n_0_0_328));
   INV_X1 i_0_0_480 (.A(n_0_0_276), .ZN(n_0_0_330));
   OAI211_X1 i_0_0_481 (.A(n_0_0_286), .B(n_0_0_331), .C1(n_0_0_338), .C2(
      n_0_0_333), .ZN(res[22]));
   AOI22_X1 i_0_0_482 (.A1(mult_res[45]), .A2(n_0_0_234), .B1(mult_res[46]), 
      .B2(n_0_0_233), .ZN(n_0_0_331));
   AOI22_X1 i_0_0_483 (.A1(mult_res[46]), .A2(n_0_0_275), .B1(mult_res[45]), 
      .B2(n_0_0_344), .ZN(n_0_0_333));
   INV_X1 i_0_0_484 (.A(n_0_0_338), .ZN(n_0_0_334));
   NAND2_X1 i_0_0_485 (.A1(n_0_0_330), .A2(n_0_0_341), .ZN(n_0_0_338));
   NOR3_X1 i_0_0_486 (.A1(n_0_0_222), .A2(n_0_0_225), .A3(n_0_0_220), .ZN(
      n_0_0_341));
   INV_X1 i_0_0_487 (.A(n_0_0_227), .ZN(n_0_0_344));
   INV_X1 i_0_0_488 (.A(mult_res[45]), .ZN(n_0_0_347));
   INV_X1 i_0_0_489 (.A(n_0_0_286), .ZN(n_0_0_370));
   OAI21_X1 i_0_0_490 (.A(n_0_0_373), .B1(n_0_0_295), .B2(n_0_0_374), .ZN(
      res[31]));
   NAND2_X1 i_0_0_491 (.A1(n_0_0_295), .A2(special_res[31]), .ZN(n_0_0_373));
   XNOR2_X1 i_0_0_492 (.A(Sa), .B(Sb), .ZN(n_0_0_374));
   AOI221_X1 i_0_0_493 (.A(n_0_0_382), .B1(n_0_0_390), .B2(n_0_0_377), .C1(
      shamt[0]), .C2(n_0_0_380), .ZN(Nb[1]));
   OAI22_X1 i_0_0_494 (.A1(n_0_59), .A2(n_0_0_73), .B1(n_0_28), .B2(n_0_0_63), 
      .ZN(n_0_0_377));
   OAI22_X1 i_0_0_495 (.A1(n_0_60), .A2(n_0_0_73), .B1(n_0_29), .B2(n_0_0_63), 
      .ZN(n_0_0_380));
   NAND2_X1 i_0_0_496 (.A1(n_0_0_393), .A2(n_0_0_386), .ZN(n_0_0_382));
   NOR3_X1 i_0_0_497 (.A1(shamt[4]), .A2(shamt[2]), .A3(shamt[3]), .ZN(n_0_0_386));
   INV_X1 i_0_0_498 (.A(shamt[0]), .ZN(n_0_0_390));
   INV_X1 i_0_0_499 (.A(shamt[1]), .ZN(n_0_0_393));
   OAI21_X1 i_0_0_500 (.A(n_0_0_396), .B1(shamt[0]), .B2(n_0_0_398), .ZN(Nb[10]));
   NAND2_X1 i_0_0_501 (.A1(shamt[0]), .A2(n_0_0_409), .ZN(n_0_0_396));
   AOI22_X1 i_0_0_502 (.A1(n_0_0_393), .A2(n_0_0_400), .B1(shamt[1]), .B2(
      n_0_0_404), .ZN(n_0_0_398));
   OAI22_X1 i_0_0_503 (.A1(n_0_0_423), .A2(n_0_0_418), .B1(shamt[2]), .B2(
      n_0_0_402), .ZN(n_0_0_400));
   AOI22_X1 i_0_0_504 (.A1(n_0_72), .A2(n_0_0_414), .B1(n_0_0_425), .B2(n_0_80), 
      .ZN(n_0_0_402));
   OAI22_X1 i_0_0_505 (.A1(n_0_0_423), .A2(n_0_0_417), .B1(shamt[2]), .B2(
      n_0_0_407), .ZN(n_0_0_404));
   AOI22_X1 i_0_0_506 (.A1(n_0_70), .A2(n_0_0_414), .B1(n_0_0_425), .B2(n_0_78), 
      .ZN(n_0_0_407));
   AOI22_X1 i_0_0_507 (.A1(n_0_0_427), .A2(n_0_0_410), .B1(n_0_0_393), .B2(
      n_0_0_411), .ZN(n_0_0_409));
   AOI22_X1 i_0_0_508 (.A1(n_0_0_386), .A2(n_0_77), .B1(n_0_0_424), .B2(n_0_73), 
      .ZN(n_0_0_410));
   INV_X1 i_0_0_509 (.A(n_0_0_412), .ZN(n_0_0_411));
   OAI22_X1 i_0_0_510 (.A1(n_0_0_426), .A2(n_0_0_423), .B1(shamt[2]), .B2(
      n_0_0_413), .ZN(n_0_0_412));
   AOI22_X1 i_0_0_511 (.A1(n_0_71), .A2(n_0_0_414), .B1(n_0_0_425), .B2(n_0_79), 
      .ZN(n_0_0_413));
   AND2_X1 i_0_0_512 (.A1(n_0_0_428), .A2(shamt[3]), .ZN(n_0_0_414));
   INV_X1 i_0_0_513 (.A(n_0_0_415), .ZN(n_0_72));
   OAI22_X1 i_0_0_514 (.A1(n_0_27), .A2(n_0_0_63), .B1(n_0_58), .B2(n_0_0_73), 
      .ZN(n_0_0_415));
   INV_X1 i_0_0_515 (.A(n_0_0_416), .ZN(n_0_73));
   OAI22_X1 i_0_0_516 (.A1(n_0_26), .A2(n_0_0_63), .B1(n_0_57), .B2(n_0_0_73), 
      .ZN(n_0_0_416));
   INV_X1 i_0_0_517 (.A(n_0_0_417), .ZN(n_0_74));
   OAI22_X1 i_0_0_518 (.A1(n_0_25), .A2(n_0_0_63), .B1(n_0_56), .B2(n_0_0_73), 
      .ZN(n_0_0_417));
   INV_X1 i_0_0_519 (.A(n_0_0_418), .ZN(n_0_76));
   OAI22_X1 i_0_0_520 (.A1(n_0_23), .A2(n_0_0_63), .B1(n_0_54), .B2(n_0_0_73), 
      .ZN(n_0_0_418));
   INV_X1 i_0_0_521 (.A(n_0_0_419), .ZN(n_0_77));
   OAI22_X1 i_0_0_522 (.A1(n_0_22), .A2(n_0_0_63), .B1(n_0_53), .B2(n_0_0_73), 
      .ZN(n_0_0_419));
   INV_X1 i_0_0_523 (.A(n_0_0_420), .ZN(n_0_78));
   AOI22_X1 i_0_0_524 (.A1(n_0_52), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_21), 
      .ZN(n_0_0_420));
   INV_X1 i_0_0_525 (.A(n_0_0_421), .ZN(n_0_79));
   AOI22_X1 i_0_0_526 (.A1(n_0_51), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_20), 
      .ZN(n_0_0_421));
   INV_X1 i_0_0_527 (.A(n_0_0_422), .ZN(n_0_80));
   AOI22_X1 i_0_0_528 (.A1(n_0_50), .A2(n_0_0_63), .B1(n_0_0_73), .B2(n_0_19), 
      .ZN(n_0_0_422));
   INV_X1 i_0_0_529 (.A(n_0_0_424), .ZN(n_0_0_423));
   NOR3_X1 i_0_0_530 (.A1(shamt[4]), .A2(shamt[3]), .A3(n_0_0_100), .ZN(
      n_0_0_424));
   NOR2_X1 i_0_0_531 (.A1(shamt[4]), .A2(shamt[3]), .ZN(n_0_0_425));
   INV_X1 i_0_0_532 (.A(n_0_0_426), .ZN(n_0_75));
   OAI22_X1 i_0_0_533 (.A1(n_0_24), .A2(n_0_0_63), .B1(n_0_55), .B2(n_0_0_73), 
      .ZN(n_0_0_426));
   INV_X1 i_0_0_534 (.A(n_0_0_380), .ZN(n_0_70));
   INV_X1 i_0_0_535 (.A(n_0_0_393), .ZN(n_0_0_427));
   INV_X1 i_0_0_536 (.A(n_0_0_377), .ZN(n_0_71));
   INV_X1 i_0_0_537 (.A(shamt[4]), .ZN(n_0_0_428));
endmodule
