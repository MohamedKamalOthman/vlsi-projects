/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 17 13:40:06 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 825441627 */

/* blackbox module registerNbits_bbox_0 */

/* blackbox module registerNbits_bbox_1 */

/* blackbox module registerNbits_bbox */

module datapath(multiplicand2, p_0);
   input [31:0]multiplicand2;
   output [31:0]p_0;

   INV_X1 i_0 (.A(multiplicand2[0]), .ZN(n_0));
   XNOR2_X1 i_1 (.A(multiplicand2[1]), .B(n_0), .ZN(p_0[1]));
   NOR2_X1 i_2 (.A1(multiplicand2[1]), .A2(multiplicand2[0]), .ZN(n_1));
   XNOR2_X1 i_3 (.A(multiplicand2[2]), .B(n_1), .ZN(p_0[2]));
   NOR2_X1 i_4 (.A1(multiplicand2[2]), .A2(n_3), .ZN(n_2));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   XNOR2_X1 i_6 (.A(multiplicand2[3]), .B(n_2), .ZN(p_0[3]));
   NOR2_X1 i_7 (.A1(multiplicand2[3]), .A2(n_5), .ZN(n_4));
   INV_X1 i_8 (.A(n_2), .ZN(n_5));
   XNOR2_X1 i_9 (.A(multiplicand2[4]), .B(n_4), .ZN(p_0[4]));
   NOR2_X1 i_10 (.A1(multiplicand2[4]), .A2(n_7), .ZN(n_6));
   INV_X1 i_11 (.A(n_4), .ZN(n_7));
   XNOR2_X1 i_12 (.A(multiplicand2[5]), .B(n_6), .ZN(p_0[5]));
   NOR2_X1 i_13 (.A1(multiplicand2[5]), .A2(n_9), .ZN(n_8));
   INV_X1 i_14 (.A(n_6), .ZN(n_9));
   XNOR2_X1 i_15 (.A(multiplicand2[6]), .B(n_8), .ZN(p_0[6]));
   NOR2_X1 i_16 (.A1(multiplicand2[6]), .A2(n_11), .ZN(n_10));
   INV_X1 i_17 (.A(n_8), .ZN(n_11));
   XNOR2_X1 i_18 (.A(multiplicand2[7]), .B(n_10), .ZN(p_0[7]));
   NOR2_X1 i_19 (.A1(multiplicand2[7]), .A2(n_13), .ZN(n_12));
   INV_X1 i_20 (.A(n_10), .ZN(n_13));
   XNOR2_X1 i_21 (.A(multiplicand2[8]), .B(n_12), .ZN(p_0[8]));
   NOR2_X1 i_22 (.A1(multiplicand2[8]), .A2(n_15), .ZN(n_14));
   INV_X1 i_23 (.A(n_12), .ZN(n_15));
   XNOR2_X1 i_24 (.A(multiplicand2[9]), .B(n_14), .ZN(p_0[9]));
   NOR2_X1 i_25 (.A1(multiplicand2[9]), .A2(n_17), .ZN(n_16));
   INV_X1 i_26 (.A(n_14), .ZN(n_17));
   XNOR2_X1 i_27 (.A(multiplicand2[10]), .B(n_16), .ZN(p_0[10]));
   NOR2_X1 i_28 (.A1(multiplicand2[10]), .A2(n_19), .ZN(n_18));
   INV_X1 i_29 (.A(n_16), .ZN(n_19));
   XNOR2_X1 i_30 (.A(multiplicand2[11]), .B(n_18), .ZN(p_0[11]));
   NOR2_X1 i_31 (.A1(multiplicand2[11]), .A2(n_21), .ZN(n_20));
   INV_X1 i_32 (.A(n_18), .ZN(n_21));
   XNOR2_X1 i_33 (.A(multiplicand2[12]), .B(n_20), .ZN(p_0[12]));
   NOR2_X1 i_34 (.A1(multiplicand2[12]), .A2(n_23), .ZN(n_22));
   INV_X1 i_35 (.A(n_20), .ZN(n_23));
   XNOR2_X1 i_36 (.A(multiplicand2[13]), .B(n_22), .ZN(p_0[13]));
   NOR2_X1 i_37 (.A1(multiplicand2[13]), .A2(n_25), .ZN(n_24));
   INV_X1 i_38 (.A(n_22), .ZN(n_25));
   XNOR2_X1 i_39 (.A(multiplicand2[14]), .B(n_24), .ZN(p_0[14]));
   NOR2_X1 i_40 (.A1(multiplicand2[14]), .A2(n_27), .ZN(n_26));
   INV_X1 i_41 (.A(n_24), .ZN(n_27));
   XNOR2_X1 i_42 (.A(multiplicand2[15]), .B(n_26), .ZN(p_0[15]));
   NOR2_X1 i_43 (.A1(multiplicand2[15]), .A2(n_29), .ZN(n_28));
   INV_X1 i_44 (.A(n_26), .ZN(n_29));
   XNOR2_X1 i_45 (.A(multiplicand2[16]), .B(n_28), .ZN(p_0[16]));
   NOR2_X1 i_46 (.A1(multiplicand2[16]), .A2(n_31), .ZN(n_30));
   INV_X1 i_47 (.A(n_28), .ZN(n_31));
   XNOR2_X1 i_48 (.A(multiplicand2[17]), .B(n_30), .ZN(p_0[17]));
   NOR2_X1 i_49 (.A1(multiplicand2[17]), .A2(n_33), .ZN(n_32));
   INV_X1 i_50 (.A(n_30), .ZN(n_33));
   XNOR2_X1 i_51 (.A(multiplicand2[18]), .B(n_32), .ZN(p_0[18]));
   NOR2_X1 i_52 (.A1(multiplicand2[18]), .A2(n_35), .ZN(n_34));
   INV_X1 i_53 (.A(n_32), .ZN(n_35));
   XNOR2_X1 i_54 (.A(multiplicand2[19]), .B(n_34), .ZN(p_0[19]));
   NOR2_X1 i_55 (.A1(multiplicand2[19]), .A2(n_37), .ZN(n_36));
   INV_X1 i_56 (.A(n_34), .ZN(n_37));
   XNOR2_X1 i_57 (.A(multiplicand2[20]), .B(n_36), .ZN(p_0[20]));
   NOR2_X1 i_58 (.A1(multiplicand2[20]), .A2(n_39), .ZN(n_38));
   INV_X1 i_59 (.A(n_36), .ZN(n_39));
   XNOR2_X1 i_60 (.A(multiplicand2[21]), .B(n_38), .ZN(p_0[21]));
   NOR2_X1 i_61 (.A1(multiplicand2[21]), .A2(n_41), .ZN(n_40));
   INV_X1 i_62 (.A(n_38), .ZN(n_41));
   XNOR2_X1 i_63 (.A(multiplicand2[22]), .B(n_40), .ZN(p_0[22]));
   NOR2_X1 i_64 (.A1(multiplicand2[22]), .A2(n_43), .ZN(n_42));
   INV_X1 i_65 (.A(n_40), .ZN(n_43));
   XNOR2_X1 i_66 (.A(multiplicand2[23]), .B(n_42), .ZN(p_0[23]));
   NOR2_X1 i_67 (.A1(multiplicand2[23]), .A2(n_45), .ZN(n_44));
   INV_X1 i_68 (.A(n_42), .ZN(n_45));
   XNOR2_X1 i_69 (.A(multiplicand2[24]), .B(n_44), .ZN(p_0[24]));
   NOR2_X1 i_70 (.A1(multiplicand2[24]), .A2(n_47), .ZN(n_46));
   INV_X1 i_71 (.A(n_44), .ZN(n_47));
   XNOR2_X1 i_72 (.A(multiplicand2[25]), .B(n_46), .ZN(p_0[25]));
   NOR2_X1 i_73 (.A1(multiplicand2[25]), .A2(n_49), .ZN(n_48));
   INV_X1 i_74 (.A(n_46), .ZN(n_49));
   XNOR2_X1 i_75 (.A(multiplicand2[26]), .B(n_48), .ZN(p_0[26]));
   NOR2_X1 i_76 (.A1(multiplicand2[26]), .A2(n_51), .ZN(n_50));
   INV_X1 i_77 (.A(n_48), .ZN(n_51));
   XNOR2_X1 i_78 (.A(multiplicand2[27]), .B(n_50), .ZN(p_0[27]));
   NOR2_X1 i_79 (.A1(multiplicand2[27]), .A2(n_53), .ZN(n_52));
   INV_X1 i_80 (.A(n_50), .ZN(n_53));
   XNOR2_X1 i_81 (.A(multiplicand2[28]), .B(n_52), .ZN(p_0[28]));
   NOR2_X1 i_82 (.A1(multiplicand2[28]), .A2(n_55), .ZN(n_54));
   INV_X1 i_83 (.A(n_52), .ZN(n_55));
   XNOR2_X1 i_84 (.A(multiplicand2[29]), .B(n_54), .ZN(p_0[29]));
   NOR2_X1 i_85 (.A1(multiplicand2[29]), .A2(n_57), .ZN(n_56));
   INV_X1 i_86 (.A(n_54), .ZN(n_57));
   XNOR2_X1 i_87 (.A(multiplicand2[30]), .B(n_56), .ZN(p_0[30]));
   NOR2_X1 i_88 (.A1(multiplicand2[30]), .A2(n_59), .ZN(n_58));
   INV_X1 i_89 (.A(n_56), .ZN(n_59));
   XNOR2_X1 i_90 (.A(multiplicand2[31]), .B(n_58), .ZN(p_0[31]));
endmodule

module datapath__0_0(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_1(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_4(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_5(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_8(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_9(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_12(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_13(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_16(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_17(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_20(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_21(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_24(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_25(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_28(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_29(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_32(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_33(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_36(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_37(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_40(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_41(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_44(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_45(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_48(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_49(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_52(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_53(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_56(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_57(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_60(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_61(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_64(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_65(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_68(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_69(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_72(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_73(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_76(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_77(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_80(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_81(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_84(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_85(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_88(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_89(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_92(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_93(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_96(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_97(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_100(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_101(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_104(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_105(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_108(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_109(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_112(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_113(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_116(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_117(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module datapath__0_120(p_0, p_1, p_2);
   input [31:0]p_0;
   input [31:0]p_1;
   output [31:0]p_2;

   INV_X1 i_0 (.A(p_0[30]), .ZN(n_0));
   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   FA_X1 i_15 (.A(p_0[14]), .B(p_1[14]), .CI(n_14), .CO(n_15), .S(p_2[14]));
   FA_X1 i_16 (.A(p_0[15]), .B(p_1[15]), .CI(n_15), .CO(n_16), .S(p_2[15]));
   FA_X1 i_17 (.A(p_0[16]), .B(p_1[16]), .CI(n_16), .CO(n_17), .S(p_2[16]));
   FA_X1 i_18 (.A(p_0[17]), .B(p_1[17]), .CI(n_17), .CO(n_18), .S(p_2[17]));
   FA_X1 i_19 (.A(p_0[18]), .B(p_1[18]), .CI(n_18), .CO(n_19), .S(p_2[18]));
   FA_X1 i_20 (.A(p_0[19]), .B(p_1[19]), .CI(n_19), .CO(n_20), .S(p_2[19]));
   FA_X1 i_21 (.A(p_0[20]), .B(p_1[20]), .CI(n_20), .CO(n_21), .S(p_2[20]));
   FA_X1 i_22 (.A(p_0[21]), .B(p_1[21]), .CI(n_21), .CO(n_22), .S(p_2[21]));
   FA_X1 i_23 (.A(p_0[22]), .B(p_1[22]), .CI(n_22), .CO(n_23), .S(p_2[22]));
   FA_X1 i_24 (.A(p_0[23]), .B(p_1[23]), .CI(n_23), .CO(n_24), .S(p_2[23]));
   FA_X1 i_25 (.A(p_0[24]), .B(p_1[24]), .CI(n_24), .CO(n_25), .S(p_2[24]));
   FA_X1 i_26 (.A(p_0[25]), .B(p_1[25]), .CI(n_25), .CO(n_26), .S(p_2[25]));
   FA_X1 i_27 (.A(p_0[26]), .B(p_1[26]), .CI(n_26), .CO(n_27), .S(p_2[26]));
   FA_X1 i_28 (.A(p_0[27]), .B(p_1[27]), .CI(n_27), .CO(n_28), .S(p_2[27]));
   FA_X1 i_29 (.A(p_0[28]), .B(p_1[28]), .CI(n_28), .CO(n_29), .S(p_2[28]));
   FA_X1 i_30 (.A(p_0[29]), .B(p_1[29]), .CI(n_29), .CO(n_30), .S(p_2[29]));
   XNOR2_X1 i_31 (.A(p_1[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_2[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_1[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(p_0[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_2[31]));
endmodule

module datapath__0_121(multiplicand2, p_0, p_1);
   input [31:0]multiplicand2;
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(multiplicand2[30]), .ZN(n_0));
   HA_X1 i_1 (.A(multiplicand2[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(multiplicand2[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(multiplicand2[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(multiplicand2[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(multiplicand2[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(multiplicand2[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(multiplicand2[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(multiplicand2[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(multiplicand2[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(multiplicand2[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(multiplicand2[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), 
      .S(p_1[10]));
   FA_X1 i_12 (.A(multiplicand2[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), 
      .S(p_1[11]));
   FA_X1 i_13 (.A(multiplicand2[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), 
      .S(p_1[12]));
   FA_X1 i_14 (.A(multiplicand2[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), 
      .S(p_1[13]));
   FA_X1 i_15 (.A(multiplicand2[14]), .B(p_0[14]), .CI(n_14), .CO(n_15), 
      .S(p_1[14]));
   FA_X1 i_16 (.A(multiplicand2[15]), .B(p_0[15]), .CI(n_15), .CO(n_16), 
      .S(p_1[15]));
   FA_X1 i_17 (.A(multiplicand2[16]), .B(p_0[16]), .CI(n_16), .CO(n_17), 
      .S(p_1[16]));
   FA_X1 i_18 (.A(multiplicand2[17]), .B(p_0[17]), .CI(n_17), .CO(n_18), 
      .S(p_1[17]));
   FA_X1 i_19 (.A(multiplicand2[18]), .B(p_0[18]), .CI(n_18), .CO(n_19), 
      .S(p_1[18]));
   FA_X1 i_20 (.A(multiplicand2[19]), .B(p_0[19]), .CI(n_19), .CO(n_20), 
      .S(p_1[19]));
   FA_X1 i_21 (.A(multiplicand2[20]), .B(p_0[20]), .CI(n_20), .CO(n_21), 
      .S(p_1[20]));
   FA_X1 i_22 (.A(multiplicand2[21]), .B(p_0[21]), .CI(n_21), .CO(n_22), 
      .S(p_1[21]));
   FA_X1 i_23 (.A(multiplicand2[22]), .B(p_0[22]), .CI(n_22), .CO(n_23), 
      .S(p_1[22]));
   FA_X1 i_24 (.A(multiplicand2[23]), .B(p_0[23]), .CI(n_23), .CO(n_24), 
      .S(p_1[23]));
   FA_X1 i_25 (.A(multiplicand2[24]), .B(p_0[24]), .CI(n_24), .CO(n_25), 
      .S(p_1[24]));
   FA_X1 i_26 (.A(multiplicand2[25]), .B(p_0[25]), .CI(n_25), .CO(n_26), 
      .S(p_1[25]));
   FA_X1 i_27 (.A(multiplicand2[26]), .B(p_0[26]), .CI(n_26), .CO(n_27), 
      .S(p_1[26]));
   FA_X1 i_28 (.A(multiplicand2[27]), .B(p_0[27]), .CI(n_27), .CO(n_28), 
      .S(p_1[27]));
   FA_X1 i_29 (.A(multiplicand2[28]), .B(p_0[28]), .CI(n_28), .CO(n_29), 
      .S(p_1[28]));
   FA_X1 i_30 (.A(multiplicand2[29]), .B(p_0[29]), .CI(n_29), .CO(n_30), 
      .S(p_1[29]));
   XNOR2_X1 i_31 (.A(p_0[30]), .B(n_0), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(n_32));
   INV_X1 i_33 (.A(n_32), .ZN(p_1[30]));
   NAND3_X1 i_34 (.A1(n_34), .A2(n_36), .A3(n_37), .ZN(n_33));
   NAND2_X1 i_35 (.A1(n_0), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(p_0[30]), .ZN(n_35));
   NAND2_X1 i_37 (.A1(n_30), .A2(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_30), .A2(n_0), .ZN(n_37));
   XNOR2_X1 i_39 (.A(multiplicand2[31]), .B(n_0), .ZN(n_38));
   XNOR2_X1 i_40 (.A(n_38), .B(n_33), .ZN(p_1[31]));
endmodule

module booth(multiplicand2, multiplier2, product);
   input [31:0]multiplicand2;
   input [31:0]multiplier2;
   output [63:0]product;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire [31:0]accumlator;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_4_0;
   wire n_0_96;
   wire n_0_97;
   wire n_0_95;
   wire n_0_5_0;
   wire n_0_5_1;
   wire n_0_98;
   wire n_0_5_2;
   wire n_0_99;
   wire n_0_5_3;
   wire n_0_100;
   wire n_0_5_4;
   wire n_0_101;
   wire n_0_5_5;
   wire n_0_102;
   wire n_0_5_6;
   wire n_0_103;
   wire n_0_5_7;
   wire n_0_104;
   wire n_0_5_8;
   wire n_0_105;
   wire n_0_5_9;
   wire n_0_106;
   wire n_0_5_10;
   wire n_0_107;
   wire n_0_5_11;
   wire n_0_108;
   wire n_0_5_12;
   wire n_0_109;
   wire n_0_5_13;
   wire n_0_110;
   wire n_0_5_14;
   wire n_0_111;
   wire n_0_5_15;
   wire n_0_112;
   wire n_0_5_16;
   wire n_0_113;
   wire n_0_5_17;
   wire n_0_114;
   wire n_0_5_18;
   wire n_0_115;
   wire n_0_5_19;
   wire n_0_116;
   wire n_0_5_20;
   wire n_0_117;
   wire n_0_5_21;
   wire n_0_118;
   wire n_0_5_22;
   wire n_0_119;
   wire n_0_5_23;
   wire n_0_120;
   wire n_0_5_24;
   wire n_0_121;
   wire n_0_5_25;
   wire n_0_122;
   wire n_0_5_26;
   wire n_0_123;
   wire n_0_5_27;
   wire n_0_124;
   wire n_0_5_28;
   wire n_0_125;
   wire n_0_5_29;
   wire n_0_126;
   wire n_0_5_30;
   wire n_0_5_31;
   wire n_0_127;
   wire n_0_5_32;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_8_0;
   wire n_0_194;
   wire n_0_195;
   wire n_0_193;
   wire n_0_9_0;
   wire n_0_9_1;
   wire n_0_196;
   wire n_0_9_2;
   wire n_0_197;
   wire n_0_9_3;
   wire n_0_198;
   wire n_0_9_4;
   wire n_0_199;
   wire n_0_9_5;
   wire n_0_200;
   wire n_0_9_6;
   wire n_0_201;
   wire n_0_9_7;
   wire n_0_202;
   wire n_0_9_8;
   wire n_0_203;
   wire n_0_9_9;
   wire n_0_204;
   wire n_0_9_10;
   wire n_0_205;
   wire n_0_9_11;
   wire n_0_206;
   wire n_0_9_12;
   wire n_0_207;
   wire n_0_9_13;
   wire n_0_208;
   wire n_0_9_14;
   wire n_0_209;
   wire n_0_9_15;
   wire n_0_210;
   wire n_0_9_16;
   wire n_0_211;
   wire n_0_9_17;
   wire n_0_212;
   wire n_0_9_18;
   wire n_0_213;
   wire n_0_9_19;
   wire n_0_214;
   wire n_0_9_20;
   wire n_0_215;
   wire n_0_9_21;
   wire n_0_216;
   wire n_0_9_22;
   wire n_0_217;
   wire n_0_9_23;
   wire n_0_218;
   wire n_0_9_24;
   wire n_0_219;
   wire n_0_9_25;
   wire n_0_220;
   wire n_0_9_26;
   wire n_0_221;
   wire n_0_9_27;
   wire n_0_222;
   wire n_0_9_28;
   wire n_0_223;
   wire n_0_9_29;
   wire n_0_224;
   wire n_0_9_30;
   wire n_0_9_31;
   wire n_0_225;
   wire n_0_9_32;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_12_0;
   wire n_0_292;
   wire n_0_293;
   wire n_0_291;
   wire n_0_13_0;
   wire n_0_13_1;
   wire n_0_294;
   wire n_0_13_2;
   wire n_0_295;
   wire n_0_13_3;
   wire n_0_296;
   wire n_0_13_4;
   wire n_0_297;
   wire n_0_13_5;
   wire n_0_298;
   wire n_0_13_6;
   wire n_0_299;
   wire n_0_13_7;
   wire n_0_300;
   wire n_0_13_8;
   wire n_0_301;
   wire n_0_13_9;
   wire n_0_302;
   wire n_0_13_10;
   wire n_0_303;
   wire n_0_13_11;
   wire n_0_304;
   wire n_0_13_12;
   wire n_0_305;
   wire n_0_13_13;
   wire n_0_306;
   wire n_0_13_14;
   wire n_0_307;
   wire n_0_13_15;
   wire n_0_308;
   wire n_0_13_16;
   wire n_0_309;
   wire n_0_13_17;
   wire n_0_310;
   wire n_0_13_18;
   wire n_0_311;
   wire n_0_13_19;
   wire n_0_312;
   wire n_0_13_20;
   wire n_0_313;
   wire n_0_13_21;
   wire n_0_314;
   wire n_0_13_22;
   wire n_0_315;
   wire n_0_13_23;
   wire n_0_316;
   wire n_0_13_24;
   wire n_0_317;
   wire n_0_13_25;
   wire n_0_318;
   wire n_0_13_26;
   wire n_0_319;
   wire n_0_13_27;
   wire n_0_320;
   wire n_0_13_28;
   wire n_0_321;
   wire n_0_13_29;
   wire n_0_322;
   wire n_0_13_30;
   wire n_0_13_31;
   wire n_0_323;
   wire n_0_13_32;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_16_0;
   wire n_0_390;
   wire n_0_391;
   wire n_0_389;
   wire n_0_17_0;
   wire n_0_17_1;
   wire n_0_392;
   wire n_0_17_2;
   wire n_0_393;
   wire n_0_17_3;
   wire n_0_394;
   wire n_0_17_4;
   wire n_0_395;
   wire n_0_17_5;
   wire n_0_396;
   wire n_0_17_6;
   wire n_0_397;
   wire n_0_17_7;
   wire n_0_398;
   wire n_0_17_8;
   wire n_0_399;
   wire n_0_17_9;
   wire n_0_400;
   wire n_0_17_10;
   wire n_0_401;
   wire n_0_17_11;
   wire n_0_402;
   wire n_0_17_12;
   wire n_0_403;
   wire n_0_17_13;
   wire n_0_404;
   wire n_0_17_14;
   wire n_0_405;
   wire n_0_17_15;
   wire n_0_406;
   wire n_0_17_16;
   wire n_0_407;
   wire n_0_17_17;
   wire n_0_408;
   wire n_0_17_18;
   wire n_0_409;
   wire n_0_17_19;
   wire n_0_410;
   wire n_0_17_20;
   wire n_0_411;
   wire n_0_17_21;
   wire n_0_412;
   wire n_0_17_22;
   wire n_0_413;
   wire n_0_17_23;
   wire n_0_414;
   wire n_0_17_24;
   wire n_0_415;
   wire n_0_17_25;
   wire n_0_416;
   wire n_0_17_26;
   wire n_0_417;
   wire n_0_17_27;
   wire n_0_418;
   wire n_0_17_28;
   wire n_0_419;
   wire n_0_17_29;
   wire n_0_420;
   wire n_0_17_30;
   wire n_0_17_31;
   wire n_0_421;
   wire n_0_17_32;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_20_0;
   wire n_0_488;
   wire n_0_489;
   wire n_0_487;
   wire n_0_21_0;
   wire n_0_21_1;
   wire n_0_490;
   wire n_0_21_2;
   wire n_0_491;
   wire n_0_21_3;
   wire n_0_492;
   wire n_0_21_4;
   wire n_0_493;
   wire n_0_21_5;
   wire n_0_494;
   wire n_0_21_6;
   wire n_0_495;
   wire n_0_21_7;
   wire n_0_496;
   wire n_0_21_8;
   wire n_0_497;
   wire n_0_21_9;
   wire n_0_498;
   wire n_0_21_10;
   wire n_0_499;
   wire n_0_21_11;
   wire n_0_500;
   wire n_0_21_12;
   wire n_0_501;
   wire n_0_21_13;
   wire n_0_502;
   wire n_0_21_14;
   wire n_0_503;
   wire n_0_21_15;
   wire n_0_504;
   wire n_0_21_16;
   wire n_0_505;
   wire n_0_21_17;
   wire n_0_506;
   wire n_0_21_18;
   wire n_0_507;
   wire n_0_21_19;
   wire n_0_508;
   wire n_0_21_20;
   wire n_0_509;
   wire n_0_21_21;
   wire n_0_510;
   wire n_0_21_22;
   wire n_0_511;
   wire n_0_21_23;
   wire n_0_512;
   wire n_0_21_24;
   wire n_0_513;
   wire n_0_21_25;
   wire n_0_514;
   wire n_0_21_26;
   wire n_0_515;
   wire n_0_21_27;
   wire n_0_516;
   wire n_0_21_28;
   wire n_0_517;
   wire n_0_21_29;
   wire n_0_518;
   wire n_0_21_30;
   wire n_0_21_31;
   wire n_0_519;
   wire n_0_21_32;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_525;
   wire n_0_526;
   wire n_0_527;
   wire n_0_528;
   wire n_0_529;
   wire n_0_530;
   wire n_0_531;
   wire n_0_532;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;
   wire n_0_537;
   wire n_0_538;
   wire n_0_539;
   wire n_0_540;
   wire n_0_541;
   wire n_0_542;
   wire n_0_543;
   wire n_0_544;
   wire n_0_545;
   wire n_0_546;
   wire n_0_547;
   wire n_0_548;
   wire n_0_549;
   wire n_0_550;
   wire n_0_551;
   wire n_0_552;
   wire n_0_553;
   wire n_0_554;
   wire n_0_555;
   wire n_0_556;
   wire n_0_557;
   wire n_0_558;
   wire n_0_559;
   wire n_0_560;
   wire n_0_561;
   wire n_0_562;
   wire n_0_563;
   wire n_0_564;
   wire n_0_565;
   wire n_0_566;
   wire n_0_567;
   wire n_0_568;
   wire n_0_569;
   wire n_0_570;
   wire n_0_571;
   wire n_0_572;
   wire n_0_573;
   wire n_0_574;
   wire n_0_575;
   wire n_0_576;
   wire n_0_577;
   wire n_0_578;
   wire n_0_579;
   wire n_0_580;
   wire n_0_581;
   wire n_0_582;
   wire n_0_583;
   wire n_0_584;
   wire n_0_24_0;
   wire n_0_586;
   wire n_0_587;
   wire n_0_585;
   wire n_0_25_0;
   wire n_0_25_1;
   wire n_0_588;
   wire n_0_25_2;
   wire n_0_589;
   wire n_0_25_3;
   wire n_0_590;
   wire n_0_25_4;
   wire n_0_591;
   wire n_0_25_5;
   wire n_0_592;
   wire n_0_25_6;
   wire n_0_593;
   wire n_0_25_7;
   wire n_0_594;
   wire n_0_25_8;
   wire n_0_595;
   wire n_0_25_9;
   wire n_0_596;
   wire n_0_25_10;
   wire n_0_597;
   wire n_0_25_11;
   wire n_0_598;
   wire n_0_25_12;
   wire n_0_599;
   wire n_0_25_13;
   wire n_0_600;
   wire n_0_25_14;
   wire n_0_601;
   wire n_0_25_15;
   wire n_0_602;
   wire n_0_25_16;
   wire n_0_603;
   wire n_0_25_17;
   wire n_0_604;
   wire n_0_25_18;
   wire n_0_605;
   wire n_0_25_19;
   wire n_0_606;
   wire n_0_25_20;
   wire n_0_607;
   wire n_0_25_21;
   wire n_0_608;
   wire n_0_25_22;
   wire n_0_609;
   wire n_0_25_23;
   wire n_0_610;
   wire n_0_25_24;
   wire n_0_611;
   wire n_0_25_25;
   wire n_0_612;
   wire n_0_25_26;
   wire n_0_613;
   wire n_0_25_27;
   wire n_0_614;
   wire n_0_25_28;
   wire n_0_615;
   wire n_0_25_29;
   wire n_0_616;
   wire n_0_25_30;
   wire n_0_25_31;
   wire n_0_617;
   wire n_0_25_32;
   wire n_0_618;
   wire n_0_619;
   wire n_0_620;
   wire n_0_621;
   wire n_0_622;
   wire n_0_623;
   wire n_0_624;
   wire n_0_625;
   wire n_0_626;
   wire n_0_627;
   wire n_0_628;
   wire n_0_629;
   wire n_0_630;
   wire n_0_631;
   wire n_0_632;
   wire n_0_633;
   wire n_0_634;
   wire n_0_635;
   wire n_0_636;
   wire n_0_637;
   wire n_0_638;
   wire n_0_639;
   wire n_0_640;
   wire n_0_641;
   wire n_0_642;
   wire n_0_643;
   wire n_0_644;
   wire n_0_645;
   wire n_0_646;
   wire n_0_647;
   wire n_0_648;
   wire n_0_649;
   wire n_0_650;
   wire n_0_651;
   wire n_0_652;
   wire n_0_653;
   wire n_0_654;
   wire n_0_655;
   wire n_0_656;
   wire n_0_657;
   wire n_0_658;
   wire n_0_659;
   wire n_0_660;
   wire n_0_661;
   wire n_0_662;
   wire n_0_663;
   wire n_0_664;
   wire n_0_665;
   wire n_0_666;
   wire n_0_667;
   wire n_0_668;
   wire n_0_669;
   wire n_0_670;
   wire n_0_671;
   wire n_0_672;
   wire n_0_673;
   wire n_0_674;
   wire n_0_675;
   wire n_0_676;
   wire n_0_677;
   wire n_0_678;
   wire n_0_679;
   wire n_0_680;
   wire n_0_681;
   wire n_0_682;
   wire n_0_28_0;
   wire n_0_684;
   wire n_0_685;
   wire n_0_683;
   wire n_0_29_0;
   wire n_0_29_1;
   wire n_0_686;
   wire n_0_29_2;
   wire n_0_687;
   wire n_0_29_3;
   wire n_0_688;
   wire n_0_29_4;
   wire n_0_689;
   wire n_0_29_5;
   wire n_0_690;
   wire n_0_29_6;
   wire n_0_691;
   wire n_0_29_7;
   wire n_0_692;
   wire n_0_29_8;
   wire n_0_693;
   wire n_0_29_9;
   wire n_0_694;
   wire n_0_29_10;
   wire n_0_695;
   wire n_0_29_11;
   wire n_0_696;
   wire n_0_29_12;
   wire n_0_697;
   wire n_0_29_13;
   wire n_0_698;
   wire n_0_29_14;
   wire n_0_699;
   wire n_0_29_15;
   wire n_0_700;
   wire n_0_29_16;
   wire n_0_701;
   wire n_0_29_17;
   wire n_0_702;
   wire n_0_29_18;
   wire n_0_703;
   wire n_0_29_19;
   wire n_0_704;
   wire n_0_29_20;
   wire n_0_705;
   wire n_0_29_21;
   wire n_0_706;
   wire n_0_29_22;
   wire n_0_707;
   wire n_0_29_23;
   wire n_0_708;
   wire n_0_29_24;
   wire n_0_709;
   wire n_0_29_25;
   wire n_0_710;
   wire n_0_29_26;
   wire n_0_711;
   wire n_0_29_27;
   wire n_0_712;
   wire n_0_29_28;
   wire n_0_713;
   wire n_0_29_29;
   wire n_0_714;
   wire n_0_29_30;
   wire n_0_29_31;
   wire n_0_715;
   wire n_0_29_32;
   wire n_0_716;
   wire n_0_717;
   wire n_0_718;
   wire n_0_719;
   wire n_0_720;
   wire n_0_721;
   wire n_0_722;
   wire n_0_723;
   wire n_0_724;
   wire n_0_725;
   wire n_0_726;
   wire n_0_727;
   wire n_0_728;
   wire n_0_729;
   wire n_0_730;
   wire n_0_731;
   wire n_0_732;
   wire n_0_733;
   wire n_0_734;
   wire n_0_735;
   wire n_0_736;
   wire n_0_737;
   wire n_0_738;
   wire n_0_739;
   wire n_0_740;
   wire n_0_741;
   wire n_0_742;
   wire n_0_743;
   wire n_0_744;
   wire n_0_745;
   wire n_0_746;
   wire n_0_747;
   wire n_0_748;
   wire n_0_749;
   wire n_0_750;
   wire n_0_751;
   wire n_0_752;
   wire n_0_753;
   wire n_0_754;
   wire n_0_755;
   wire n_0_756;
   wire n_0_757;
   wire n_0_758;
   wire n_0_759;
   wire n_0_760;
   wire n_0_761;
   wire n_0_762;
   wire n_0_763;
   wire n_0_764;
   wire n_0_765;
   wire n_0_766;
   wire n_0_767;
   wire n_0_768;
   wire n_0_769;
   wire n_0_770;
   wire n_0_771;
   wire n_0_772;
   wire n_0_773;
   wire n_0_774;
   wire n_0_775;
   wire n_0_776;
   wire n_0_777;
   wire n_0_778;
   wire n_0_779;
   wire n_0_780;
   wire n_0_32_0;
   wire n_0_782;
   wire n_0_783;
   wire n_0_781;
   wire n_0_33_0;
   wire n_0_33_1;
   wire n_0_784;
   wire n_0_33_2;
   wire n_0_785;
   wire n_0_33_3;
   wire n_0_786;
   wire n_0_33_4;
   wire n_0_787;
   wire n_0_33_5;
   wire n_0_788;
   wire n_0_33_6;
   wire n_0_789;
   wire n_0_33_7;
   wire n_0_790;
   wire n_0_33_8;
   wire n_0_791;
   wire n_0_33_9;
   wire n_0_792;
   wire n_0_33_10;
   wire n_0_793;
   wire n_0_33_11;
   wire n_0_794;
   wire n_0_33_12;
   wire n_0_795;
   wire n_0_33_13;
   wire n_0_796;
   wire n_0_33_14;
   wire n_0_797;
   wire n_0_33_15;
   wire n_0_798;
   wire n_0_33_16;
   wire n_0_799;
   wire n_0_33_17;
   wire n_0_800;
   wire n_0_33_18;
   wire n_0_801;
   wire n_0_33_19;
   wire n_0_802;
   wire n_0_33_20;
   wire n_0_803;
   wire n_0_33_21;
   wire n_0_804;
   wire n_0_33_22;
   wire n_0_805;
   wire n_0_33_23;
   wire n_0_806;
   wire n_0_33_24;
   wire n_0_807;
   wire n_0_33_25;
   wire n_0_808;
   wire n_0_33_26;
   wire n_0_809;
   wire n_0_33_27;
   wire n_0_810;
   wire n_0_33_28;
   wire n_0_811;
   wire n_0_33_29;
   wire n_0_812;
   wire n_0_33_30;
   wire n_0_33_31;
   wire n_0_813;
   wire n_0_33_32;
   wire n_0_814;
   wire n_0_815;
   wire n_0_816;
   wire n_0_817;
   wire n_0_818;
   wire n_0_819;
   wire n_0_820;
   wire n_0_821;
   wire n_0_822;
   wire n_0_823;
   wire n_0_824;
   wire n_0_825;
   wire n_0_826;
   wire n_0_827;
   wire n_0_828;
   wire n_0_829;
   wire n_0_830;
   wire n_0_831;
   wire n_0_832;
   wire n_0_833;
   wire n_0_834;
   wire n_0_835;
   wire n_0_836;
   wire n_0_837;
   wire n_0_838;
   wire n_0_839;
   wire n_0_840;
   wire n_0_841;
   wire n_0_842;
   wire n_0_843;
   wire n_0_844;
   wire n_0_845;
   wire n_0_846;
   wire n_0_847;
   wire n_0_848;
   wire n_0_849;
   wire n_0_850;
   wire n_0_851;
   wire n_0_852;
   wire n_0_853;
   wire n_0_854;
   wire n_0_855;
   wire n_0_856;
   wire n_0_857;
   wire n_0_858;
   wire n_0_859;
   wire n_0_860;
   wire n_0_861;
   wire n_0_862;
   wire n_0_863;
   wire n_0_864;
   wire n_0_865;
   wire n_0_866;
   wire n_0_867;
   wire n_0_868;
   wire n_0_869;
   wire n_0_870;
   wire n_0_871;
   wire n_0_872;
   wire n_0_873;
   wire n_0_874;
   wire n_0_875;
   wire n_0_876;
   wire n_0_877;
   wire n_0_878;
   wire n_0_36_0;
   wire n_0_880;
   wire n_0_881;
   wire n_0_879;
   wire n_0_37_0;
   wire n_0_37_1;
   wire n_0_882;
   wire n_0_37_2;
   wire n_0_883;
   wire n_0_37_3;
   wire n_0_884;
   wire n_0_37_4;
   wire n_0_885;
   wire n_0_37_5;
   wire n_0_886;
   wire n_0_37_6;
   wire n_0_887;
   wire n_0_37_7;
   wire n_0_888;
   wire n_0_37_8;
   wire n_0_889;
   wire n_0_37_9;
   wire n_0_890;
   wire n_0_37_10;
   wire n_0_891;
   wire n_0_37_11;
   wire n_0_892;
   wire n_0_37_12;
   wire n_0_893;
   wire n_0_37_13;
   wire n_0_894;
   wire n_0_37_14;
   wire n_0_895;
   wire n_0_37_15;
   wire n_0_896;
   wire n_0_37_16;
   wire n_0_897;
   wire n_0_37_17;
   wire n_0_898;
   wire n_0_37_18;
   wire n_0_899;
   wire n_0_37_19;
   wire n_0_900;
   wire n_0_37_20;
   wire n_0_901;
   wire n_0_37_21;
   wire n_0_902;
   wire n_0_37_22;
   wire n_0_903;
   wire n_0_37_23;
   wire n_0_904;
   wire n_0_37_24;
   wire n_0_905;
   wire n_0_37_25;
   wire n_0_906;
   wire n_0_37_26;
   wire n_0_907;
   wire n_0_37_27;
   wire n_0_908;
   wire n_0_37_28;
   wire n_0_909;
   wire n_0_37_29;
   wire n_0_910;
   wire n_0_37_30;
   wire n_0_37_31;
   wire n_0_911;
   wire n_0_37_32;
   wire n_0_912;
   wire n_0_913;
   wire n_0_914;
   wire n_0_915;
   wire n_0_916;
   wire n_0_917;
   wire n_0_918;
   wire n_0_919;
   wire n_0_920;
   wire n_0_921;
   wire n_0_922;
   wire n_0_923;
   wire n_0_924;
   wire n_0_925;
   wire n_0_926;
   wire n_0_927;
   wire n_0_928;
   wire n_0_929;
   wire n_0_930;
   wire n_0_931;
   wire n_0_932;
   wire n_0_933;
   wire n_0_934;
   wire n_0_935;
   wire n_0_936;
   wire n_0_937;
   wire n_0_938;
   wire n_0_939;
   wire n_0_940;
   wire n_0_941;
   wire n_0_942;
   wire n_0_943;
   wire n_0_944;
   wire n_0_945;
   wire n_0_946;
   wire n_0_947;
   wire n_0_948;
   wire n_0_949;
   wire n_0_950;
   wire n_0_951;
   wire n_0_952;
   wire n_0_953;
   wire n_0_954;
   wire n_0_955;
   wire n_0_956;
   wire n_0_957;
   wire n_0_958;
   wire n_0_959;
   wire n_0_960;
   wire n_0_961;
   wire n_0_962;
   wire n_0_963;
   wire n_0_964;
   wire n_0_965;
   wire n_0_966;
   wire n_0_967;
   wire n_0_968;
   wire n_0_969;
   wire n_0_970;
   wire n_0_971;
   wire n_0_972;
   wire n_0_973;
   wire n_0_974;
   wire n_0_975;
   wire n_0_976;
   wire n_0_40_0;
   wire n_0_978;
   wire n_0_979;
   wire n_0_977;
   wire n_0_41_0;
   wire n_0_41_1;
   wire n_0_980;
   wire n_0_41_2;
   wire n_0_981;
   wire n_0_41_3;
   wire n_0_982;
   wire n_0_41_4;
   wire n_0_983;
   wire n_0_41_5;
   wire n_0_984;
   wire n_0_41_6;
   wire n_0_985;
   wire n_0_41_7;
   wire n_0_986;
   wire n_0_41_8;
   wire n_0_987;
   wire n_0_41_9;
   wire n_0_988;
   wire n_0_41_10;
   wire n_0_989;
   wire n_0_41_11;
   wire n_0_990;
   wire n_0_41_12;
   wire n_0_991;
   wire n_0_41_13;
   wire n_0_992;
   wire n_0_41_14;
   wire n_0_993;
   wire n_0_41_15;
   wire n_0_994;
   wire n_0_41_16;
   wire n_0_995;
   wire n_0_41_17;
   wire n_0_996;
   wire n_0_41_18;
   wire n_0_997;
   wire n_0_41_19;
   wire n_0_998;
   wire n_0_41_20;
   wire n_0_999;
   wire n_0_41_21;
   wire n_0_1000;
   wire n_0_41_22;
   wire n_0_1001;
   wire n_0_41_23;
   wire n_0_1002;
   wire n_0_41_24;
   wire n_0_1003;
   wire n_0_41_25;
   wire n_0_1004;
   wire n_0_41_26;
   wire n_0_1005;
   wire n_0_41_27;
   wire n_0_1006;
   wire n_0_41_28;
   wire n_0_1007;
   wire n_0_41_29;
   wire n_0_1008;
   wire n_0_41_30;
   wire n_0_41_31;
   wire n_0_1009;
   wire n_0_41_32;
   wire n_0_1010;
   wire n_0_1011;
   wire n_0_1012;
   wire n_0_1013;
   wire n_0_1014;
   wire n_0_1015;
   wire n_0_1016;
   wire n_0_1017;
   wire n_0_1018;
   wire n_0_1019;
   wire n_0_1020;
   wire n_0_1021;
   wire n_0_1022;
   wire n_0_1023;
   wire n_0_1024;
   wire n_0_1025;
   wire n_0_1026;
   wire n_0_1027;
   wire n_0_1028;
   wire n_0_1029;
   wire n_0_1030;
   wire n_0_1031;
   wire n_0_1032;
   wire n_0_1033;
   wire n_0_1034;
   wire n_0_1035;
   wire n_0_1036;
   wire n_0_1037;
   wire n_0_1038;
   wire n_0_1039;
   wire n_0_1040;
   wire n_0_1041;
   wire n_0_1042;
   wire n_0_1043;
   wire n_0_1044;
   wire n_0_1045;
   wire n_0_1046;
   wire n_0_1047;
   wire n_0_1048;
   wire n_0_1049;
   wire n_0_1050;
   wire n_0_1051;
   wire n_0_1052;
   wire n_0_1053;
   wire n_0_1054;
   wire n_0_1055;
   wire n_0_1056;
   wire n_0_1057;
   wire n_0_1058;
   wire n_0_1059;
   wire n_0_1060;
   wire n_0_1061;
   wire n_0_1062;
   wire n_0_1063;
   wire n_0_1064;
   wire n_0_1065;
   wire n_0_1066;
   wire n_0_1067;
   wire n_0_1068;
   wire n_0_1069;
   wire n_0_1070;
   wire n_0_1071;
   wire n_0_1072;
   wire n_0_1073;
   wire n_0_1074;
   wire n_0_44_0;
   wire n_0_1076;
   wire n_0_1077;
   wire n_0_1075;
   wire n_0_45_0;
   wire n_0_45_1;
   wire n_0_1078;
   wire n_0_45_2;
   wire n_0_1079;
   wire n_0_45_3;
   wire n_0_1080;
   wire n_0_45_4;
   wire n_0_1081;
   wire n_0_45_5;
   wire n_0_1082;
   wire n_0_45_6;
   wire n_0_1083;
   wire n_0_45_7;
   wire n_0_1084;
   wire n_0_45_8;
   wire n_0_1085;
   wire n_0_45_9;
   wire n_0_1086;
   wire n_0_45_10;
   wire n_0_1087;
   wire n_0_45_11;
   wire n_0_1088;
   wire n_0_45_12;
   wire n_0_1089;
   wire n_0_45_13;
   wire n_0_1090;
   wire n_0_45_14;
   wire n_0_1091;
   wire n_0_45_15;
   wire n_0_1092;
   wire n_0_45_16;
   wire n_0_1093;
   wire n_0_45_17;
   wire n_0_1094;
   wire n_0_45_18;
   wire n_0_1095;
   wire n_0_45_19;
   wire n_0_1096;
   wire n_0_45_20;
   wire n_0_1097;
   wire n_0_45_21;
   wire n_0_1098;
   wire n_0_45_22;
   wire n_0_1099;
   wire n_0_45_23;
   wire n_0_1100;
   wire n_0_45_24;
   wire n_0_1101;
   wire n_0_45_25;
   wire n_0_1102;
   wire n_0_45_26;
   wire n_0_1103;
   wire n_0_45_27;
   wire n_0_1104;
   wire n_0_45_28;
   wire n_0_1105;
   wire n_0_45_29;
   wire n_0_1106;
   wire n_0_45_30;
   wire n_0_45_31;
   wire n_0_1107;
   wire n_0_45_32;
   wire n_0_1108;
   wire n_0_1109;
   wire n_0_1110;
   wire n_0_1111;
   wire n_0_1112;
   wire n_0_1113;
   wire n_0_1114;
   wire n_0_1115;
   wire n_0_1116;
   wire n_0_1117;
   wire n_0_1118;
   wire n_0_1119;
   wire n_0_1120;
   wire n_0_1121;
   wire n_0_1122;
   wire n_0_1123;
   wire n_0_1124;
   wire n_0_1125;
   wire n_0_1126;
   wire n_0_1127;
   wire n_0_1128;
   wire n_0_1129;
   wire n_0_1130;
   wire n_0_1131;
   wire n_0_1132;
   wire n_0_1133;
   wire n_0_1134;
   wire n_0_1135;
   wire n_0_1136;
   wire n_0_1137;
   wire n_0_1138;
   wire n_0_1139;
   wire n_0_1140;
   wire n_0_1141;
   wire n_0_1142;
   wire n_0_1143;
   wire n_0_1144;
   wire n_0_1145;
   wire n_0_1146;
   wire n_0_1147;
   wire n_0_1148;
   wire n_0_1149;
   wire n_0_1150;
   wire n_0_1151;
   wire n_0_1152;
   wire n_0_1153;
   wire n_0_1154;
   wire n_0_1155;
   wire n_0_1156;
   wire n_0_1157;
   wire n_0_1158;
   wire n_0_1159;
   wire n_0_1160;
   wire n_0_1161;
   wire n_0_1162;
   wire n_0_1163;
   wire n_0_1164;
   wire n_0_1165;
   wire n_0_1166;
   wire n_0_1167;
   wire n_0_1168;
   wire n_0_1169;
   wire n_0_1170;
   wire n_0_1171;
   wire n_0_1172;
   wire n_0_48_0;
   wire n_0_1174;
   wire n_0_1175;
   wire n_0_1173;
   wire n_0_49_0;
   wire n_0_49_1;
   wire n_0_1176;
   wire n_0_49_2;
   wire n_0_1177;
   wire n_0_49_3;
   wire n_0_1178;
   wire n_0_49_4;
   wire n_0_1179;
   wire n_0_49_5;
   wire n_0_1180;
   wire n_0_49_6;
   wire n_0_1181;
   wire n_0_49_7;
   wire n_0_1182;
   wire n_0_49_8;
   wire n_0_1183;
   wire n_0_49_9;
   wire n_0_1184;
   wire n_0_49_10;
   wire n_0_1185;
   wire n_0_49_11;
   wire n_0_1186;
   wire n_0_49_12;
   wire n_0_1187;
   wire n_0_49_13;
   wire n_0_1188;
   wire n_0_49_14;
   wire n_0_1189;
   wire n_0_49_15;
   wire n_0_1190;
   wire n_0_49_16;
   wire n_0_1191;
   wire n_0_49_17;
   wire n_0_1192;
   wire n_0_49_18;
   wire n_0_1193;
   wire n_0_49_19;
   wire n_0_1194;
   wire n_0_49_20;
   wire n_0_1195;
   wire n_0_49_21;
   wire n_0_1196;
   wire n_0_49_22;
   wire n_0_1197;
   wire n_0_49_23;
   wire n_0_1198;
   wire n_0_49_24;
   wire n_0_1199;
   wire n_0_49_25;
   wire n_0_1200;
   wire n_0_49_26;
   wire n_0_1201;
   wire n_0_49_27;
   wire n_0_1202;
   wire n_0_49_28;
   wire n_0_1203;
   wire n_0_49_29;
   wire n_0_1204;
   wire n_0_49_30;
   wire n_0_49_31;
   wire n_0_1205;
   wire n_0_49_32;
   wire n_0_1206;
   wire n_0_1207;
   wire n_0_1208;
   wire n_0_1209;
   wire n_0_1210;
   wire n_0_1211;
   wire n_0_1212;
   wire n_0_1213;
   wire n_0_1214;
   wire n_0_1215;
   wire n_0_1216;
   wire n_0_1217;
   wire n_0_1218;
   wire n_0_1219;
   wire n_0_1220;
   wire n_0_1221;
   wire n_0_1222;
   wire n_0_1223;
   wire n_0_1224;
   wire n_0_1225;
   wire n_0_1226;
   wire n_0_1227;
   wire n_0_1228;
   wire n_0_1229;
   wire n_0_1230;
   wire n_0_1231;
   wire n_0_1232;
   wire n_0_1233;
   wire n_0_1234;
   wire n_0_1235;
   wire n_0_1236;
   wire n_0_1237;
   wire n_0_1238;
   wire n_0_1239;
   wire n_0_1240;
   wire n_0_1241;
   wire n_0_1242;
   wire n_0_1243;
   wire n_0_1244;
   wire n_0_1245;
   wire n_0_1246;
   wire n_0_1247;
   wire n_0_1248;
   wire n_0_1249;
   wire n_0_1250;
   wire n_0_1251;
   wire n_0_1252;
   wire n_0_1253;
   wire n_0_1254;
   wire n_0_1255;
   wire n_0_1256;
   wire n_0_1257;
   wire n_0_1258;
   wire n_0_1259;
   wire n_0_1260;
   wire n_0_1261;
   wire n_0_1262;
   wire n_0_1263;
   wire n_0_1264;
   wire n_0_1265;
   wire n_0_1266;
   wire n_0_1267;
   wire n_0_1268;
   wire n_0_1269;
   wire n_0_1270;
   wire n_0_52_0;
   wire n_0_1272;
   wire n_0_1273;
   wire n_0_1271;
   wire n_0_53_0;
   wire n_0_53_1;
   wire n_0_1274;
   wire n_0_53_2;
   wire n_0_1275;
   wire n_0_53_3;
   wire n_0_1276;
   wire n_0_53_4;
   wire n_0_1277;
   wire n_0_53_5;
   wire n_0_1278;
   wire n_0_53_6;
   wire n_0_1279;
   wire n_0_53_7;
   wire n_0_1280;
   wire n_0_53_8;
   wire n_0_1281;
   wire n_0_53_9;
   wire n_0_1282;
   wire n_0_53_10;
   wire n_0_1283;
   wire n_0_53_11;
   wire n_0_1284;
   wire n_0_53_12;
   wire n_0_1285;
   wire n_0_53_13;
   wire n_0_1286;
   wire n_0_53_14;
   wire n_0_1287;
   wire n_0_53_15;
   wire n_0_1288;
   wire n_0_53_16;
   wire n_0_1289;
   wire n_0_53_17;
   wire n_0_1290;
   wire n_0_53_18;
   wire n_0_1291;
   wire n_0_53_19;
   wire n_0_1292;
   wire n_0_53_20;
   wire n_0_1293;
   wire n_0_53_21;
   wire n_0_1294;
   wire n_0_53_22;
   wire n_0_1295;
   wire n_0_53_23;
   wire n_0_1296;
   wire n_0_53_24;
   wire n_0_1297;
   wire n_0_53_25;
   wire n_0_1298;
   wire n_0_53_26;
   wire n_0_1299;
   wire n_0_53_27;
   wire n_0_1300;
   wire n_0_53_28;
   wire n_0_1301;
   wire n_0_53_29;
   wire n_0_1302;
   wire n_0_53_30;
   wire n_0_53_31;
   wire n_0_1303;
   wire n_0_53_32;
   wire n_0_1304;
   wire n_0_1305;
   wire n_0_1306;
   wire n_0_1307;
   wire n_0_1308;
   wire n_0_1309;
   wire n_0_1310;
   wire n_0_1311;
   wire n_0_1312;
   wire n_0_1313;
   wire n_0_1314;
   wire n_0_1315;
   wire n_0_1316;
   wire n_0_1317;
   wire n_0_1318;
   wire n_0_1319;
   wire n_0_1320;
   wire n_0_1321;
   wire n_0_1322;
   wire n_0_1323;
   wire n_0_1324;
   wire n_0_1325;
   wire n_0_1326;
   wire n_0_1327;
   wire n_0_1328;
   wire n_0_1329;
   wire n_0_1330;
   wire n_0_1331;
   wire n_0_1332;
   wire n_0_1333;
   wire n_0_1334;
   wire n_0_1335;
   wire n_0_1336;
   wire n_0_1337;
   wire n_0_1338;
   wire n_0_1339;
   wire n_0_1340;
   wire n_0_1341;
   wire n_0_1342;
   wire n_0_1343;
   wire n_0_1344;
   wire n_0_1345;
   wire n_0_1346;
   wire n_0_1347;
   wire n_0_1348;
   wire n_0_1349;
   wire n_0_1350;
   wire n_0_1351;
   wire n_0_1352;
   wire n_0_1353;
   wire n_0_1354;
   wire n_0_1355;
   wire n_0_1356;
   wire n_0_1357;
   wire n_0_1358;
   wire n_0_1359;
   wire n_0_1360;
   wire n_0_1361;
   wire n_0_1362;
   wire n_0_1363;
   wire n_0_1364;
   wire n_0_1365;
   wire n_0_1366;
   wire n_0_1367;
   wire n_0_1368;
   wire n_0_56_0;
   wire n_0_1370;
   wire n_0_1371;
   wire n_0_1369;
   wire n_0_57_0;
   wire n_0_57_1;
   wire n_0_1372;
   wire n_0_57_2;
   wire n_0_1373;
   wire n_0_57_3;
   wire n_0_1374;
   wire n_0_57_4;
   wire n_0_1375;
   wire n_0_57_5;
   wire n_0_1376;
   wire n_0_57_6;
   wire n_0_1377;
   wire n_0_57_7;
   wire n_0_1378;
   wire n_0_57_8;
   wire n_0_1379;
   wire n_0_57_9;
   wire n_0_1380;
   wire n_0_57_10;
   wire n_0_1381;
   wire n_0_57_11;
   wire n_0_1382;
   wire n_0_57_12;
   wire n_0_1383;
   wire n_0_57_13;
   wire n_0_1384;
   wire n_0_57_14;
   wire n_0_1385;
   wire n_0_57_15;
   wire n_0_1386;
   wire n_0_57_16;
   wire n_0_1387;
   wire n_0_57_17;
   wire n_0_1388;
   wire n_0_57_18;
   wire n_0_1389;
   wire n_0_57_19;
   wire n_0_1390;
   wire n_0_57_20;
   wire n_0_1391;
   wire n_0_57_21;
   wire n_0_1392;
   wire n_0_57_22;
   wire n_0_1393;
   wire n_0_57_23;
   wire n_0_1394;
   wire n_0_57_24;
   wire n_0_1395;
   wire n_0_57_25;
   wire n_0_1396;
   wire n_0_57_26;
   wire n_0_1397;
   wire n_0_57_27;
   wire n_0_1398;
   wire n_0_57_28;
   wire n_0_1399;
   wire n_0_57_29;
   wire n_0_1400;
   wire n_0_57_30;
   wire n_0_57_31;
   wire n_0_1401;
   wire n_0_57_32;
   wire n_0_1402;
   wire n_0_1403;
   wire n_0_1404;
   wire n_0_1405;
   wire n_0_1406;
   wire n_0_1407;
   wire n_0_1408;
   wire n_0_1409;
   wire n_0_1410;
   wire n_0_1411;
   wire n_0_1412;
   wire n_0_1413;
   wire n_0_1414;
   wire n_0_1415;
   wire n_0_1416;
   wire n_0_1417;
   wire n_0_1418;
   wire n_0_1419;
   wire n_0_1420;
   wire n_0_1421;
   wire n_0_1422;
   wire n_0_1423;
   wire n_0_1424;
   wire n_0_1425;
   wire n_0_1426;
   wire n_0_1427;
   wire n_0_1428;
   wire n_0_1429;
   wire n_0_1430;
   wire n_0_1431;
   wire n_0_1432;
   wire n_0_1433;
   wire n_0_1434;
   wire n_0_1435;
   wire n_0_1436;
   wire n_0_1437;
   wire n_0_1438;
   wire n_0_1439;
   wire n_0_1440;
   wire n_0_1441;
   wire n_0_1442;
   wire n_0_1443;
   wire n_0_1444;
   wire n_0_1445;
   wire n_0_1446;
   wire n_0_1447;
   wire n_0_1448;
   wire n_0_1449;
   wire n_0_1450;
   wire n_0_1451;
   wire n_0_1452;
   wire n_0_1453;
   wire n_0_1454;
   wire n_0_1455;
   wire n_0_1456;
   wire n_0_1457;
   wire n_0_1458;
   wire n_0_1459;
   wire n_0_1460;
   wire n_0_1461;
   wire n_0_1462;
   wire n_0_1463;
   wire n_0_1464;
   wire n_0_1465;
   wire n_0_1466;
   wire n_0_60_0;
   wire n_0_1468;
   wire n_0_1469;
   wire n_0_1467;
   wire n_0_61_0;
   wire n_0_61_1;
   wire n_0_1470;
   wire n_0_61_2;
   wire n_0_1471;
   wire n_0_61_3;
   wire n_0_1472;
   wire n_0_61_4;
   wire n_0_1473;
   wire n_0_61_5;
   wire n_0_1474;
   wire n_0_61_6;
   wire n_0_1475;
   wire n_0_61_7;
   wire n_0_1476;
   wire n_0_61_8;
   wire n_0_1477;
   wire n_0_61_9;
   wire n_0_1478;
   wire n_0_61_10;
   wire n_0_1479;
   wire n_0_61_11;
   wire n_0_1480;
   wire n_0_61_12;
   wire n_0_1481;
   wire n_0_61_13;
   wire n_0_1482;
   wire n_0_61_14;
   wire n_0_1483;
   wire n_0_61_15;
   wire n_0_1484;
   wire n_0_61_16;
   wire n_0_1485;
   wire n_0_61_17;
   wire n_0_1486;
   wire n_0_61_18;
   wire n_0_1487;
   wire n_0_61_19;
   wire n_0_1488;
   wire n_0_61_20;
   wire n_0_1489;
   wire n_0_61_21;
   wire n_0_1490;
   wire n_0_61_22;
   wire n_0_1491;
   wire n_0_61_23;
   wire n_0_1492;
   wire n_0_61_24;
   wire n_0_1493;
   wire n_0_61_25;
   wire n_0_1494;
   wire n_0_61_26;
   wire n_0_1495;
   wire n_0_61_27;
   wire n_0_1496;
   wire n_0_61_28;
   wire n_0_1497;
   wire n_0_61_29;
   wire n_0_1498;
   wire n_0_61_30;
   wire n_0_61_31;
   wire n_0_1499;
   wire n_0_61_32;
   wire n_0_1500;
   wire n_0_1501;
   wire n_0_1502;
   wire n_0_1503;
   wire n_0_1504;
   wire n_0_1505;
   wire n_0_1506;
   wire n_0_1507;
   wire n_0_1508;
   wire n_0_1509;
   wire n_0_1510;
   wire n_0_1511;
   wire n_0_1512;
   wire n_0_1513;
   wire n_0_1514;
   wire n_0_1515;
   wire n_0_1516;
   wire n_0_1517;
   wire n_0_1518;
   wire n_0_1519;
   wire n_0_1520;
   wire n_0_1521;
   wire n_0_1522;
   wire n_0_1523;
   wire n_0_1524;
   wire n_0_1525;
   wire n_0_1526;
   wire n_0_1527;
   wire n_0_1528;
   wire n_0_1529;
   wire n_0_1530;
   wire n_0_1531;
   wire n_0_1532;
   wire n_0_1533;
   wire n_0_1534;
   wire n_0_1535;
   wire n_0_1536;
   wire n_0_1537;
   wire n_0_1538;
   wire n_0_1539;
   wire n_0_1540;
   wire n_0_1541;
   wire n_0_1542;
   wire n_0_1543;
   wire n_0_1544;
   wire n_0_1545;
   wire n_0_1546;
   wire n_0_1547;
   wire n_0_1548;
   wire n_0_1549;
   wire n_0_1550;
   wire n_0_1551;
   wire n_0_1552;
   wire n_0_1553;
   wire n_0_1554;
   wire n_0_1555;
   wire n_0_1556;
   wire n_0_1557;
   wire n_0_1558;
   wire n_0_1559;
   wire n_0_1560;
   wire n_0_1561;
   wire n_0_1562;
   wire n_0_1563;
   wire n_0_1564;
   wire n_0_64_0;
   wire n_0_1566;
   wire n_0_1567;
   wire n_0_1565;
   wire n_0_65_0;
   wire n_0_65_1;
   wire n_0_1568;
   wire n_0_65_2;
   wire n_0_1569;
   wire n_0_65_3;
   wire n_0_1570;
   wire n_0_65_4;
   wire n_0_1571;
   wire n_0_65_5;
   wire n_0_1572;
   wire n_0_65_6;
   wire n_0_1573;
   wire n_0_65_7;
   wire n_0_1574;
   wire n_0_65_8;
   wire n_0_1575;
   wire n_0_65_9;
   wire n_0_1576;
   wire n_0_65_10;
   wire n_0_1577;
   wire n_0_65_11;
   wire n_0_1578;
   wire n_0_65_12;
   wire n_0_1579;
   wire n_0_65_13;
   wire n_0_1580;
   wire n_0_65_14;
   wire n_0_1581;
   wire n_0_65_15;
   wire n_0_1582;
   wire n_0_65_16;
   wire n_0_1583;
   wire n_0_65_17;
   wire n_0_1584;
   wire n_0_65_18;
   wire n_0_1585;
   wire n_0_65_19;
   wire n_0_1586;
   wire n_0_65_20;
   wire n_0_1587;
   wire n_0_65_21;
   wire n_0_1588;
   wire n_0_65_22;
   wire n_0_1589;
   wire n_0_65_23;
   wire n_0_1590;
   wire n_0_65_24;
   wire n_0_1591;
   wire n_0_65_25;
   wire n_0_1592;
   wire n_0_65_26;
   wire n_0_1593;
   wire n_0_65_27;
   wire n_0_1594;
   wire n_0_65_28;
   wire n_0_1595;
   wire n_0_65_29;
   wire n_0_1596;
   wire n_0_65_30;
   wire n_0_65_31;
   wire n_0_1597;
   wire n_0_65_32;
   wire n_0_1598;
   wire n_0_1599;
   wire n_0_1600;
   wire n_0_1601;
   wire n_0_1602;
   wire n_0_1603;
   wire n_0_1604;
   wire n_0_1605;
   wire n_0_1606;
   wire n_0_1607;
   wire n_0_1608;
   wire n_0_1609;
   wire n_0_1610;
   wire n_0_1611;
   wire n_0_1612;
   wire n_0_1613;
   wire n_0_1614;
   wire n_0_1615;
   wire n_0_1616;
   wire n_0_1617;
   wire n_0_1618;
   wire n_0_1619;
   wire n_0_1620;
   wire n_0_1621;
   wire n_0_1622;
   wire n_0_1623;
   wire n_0_1624;
   wire n_0_1625;
   wire n_0_1626;
   wire n_0_1627;
   wire n_0_1628;
   wire n_0_1629;
   wire n_0_1630;
   wire n_0_1631;
   wire n_0_1632;
   wire n_0_1633;
   wire n_0_1634;
   wire n_0_1635;
   wire n_0_1636;
   wire n_0_1637;
   wire n_0_1638;
   wire n_0_1639;
   wire n_0_1640;
   wire n_0_1641;
   wire n_0_1642;
   wire n_0_1643;
   wire n_0_1644;
   wire n_0_1645;
   wire n_0_1646;
   wire n_0_1647;
   wire n_0_1648;
   wire n_0_1649;
   wire n_0_1650;
   wire n_0_1651;
   wire n_0_1652;
   wire n_0_1653;
   wire n_0_1654;
   wire n_0_1655;
   wire n_0_1656;
   wire n_0_1657;
   wire n_0_1658;
   wire n_0_1659;
   wire n_0_1660;
   wire n_0_1661;
   wire n_0_1662;
   wire n_0_68_0;
   wire n_0_1664;
   wire n_0_1665;
   wire n_0_1663;
   wire n_0_69_0;
   wire n_0_69_1;
   wire n_0_1666;
   wire n_0_69_2;
   wire n_0_1667;
   wire n_0_69_3;
   wire n_0_1668;
   wire n_0_69_4;
   wire n_0_1669;
   wire n_0_69_5;
   wire n_0_1670;
   wire n_0_69_6;
   wire n_0_1671;
   wire n_0_69_7;
   wire n_0_1672;
   wire n_0_69_8;
   wire n_0_1673;
   wire n_0_69_9;
   wire n_0_1674;
   wire n_0_69_10;
   wire n_0_1675;
   wire n_0_69_11;
   wire n_0_1676;
   wire n_0_69_12;
   wire n_0_1677;
   wire n_0_69_13;
   wire n_0_1678;
   wire n_0_69_14;
   wire n_0_1679;
   wire n_0_69_15;
   wire n_0_1680;
   wire n_0_69_16;
   wire n_0_1681;
   wire n_0_69_17;
   wire n_0_1682;
   wire n_0_69_18;
   wire n_0_1683;
   wire n_0_69_19;
   wire n_0_1684;
   wire n_0_69_20;
   wire n_0_1685;
   wire n_0_69_21;
   wire n_0_1686;
   wire n_0_69_22;
   wire n_0_1687;
   wire n_0_69_23;
   wire n_0_1688;
   wire n_0_69_24;
   wire n_0_1689;
   wire n_0_69_25;
   wire n_0_1690;
   wire n_0_69_26;
   wire n_0_1691;
   wire n_0_69_27;
   wire n_0_1692;
   wire n_0_69_28;
   wire n_0_1693;
   wire n_0_69_29;
   wire n_0_1694;
   wire n_0_69_30;
   wire n_0_69_31;
   wire n_0_1695;
   wire n_0_69_32;
   wire n_0_1696;
   wire n_0_1697;
   wire n_0_1698;
   wire n_0_1699;
   wire n_0_1700;
   wire n_0_1701;
   wire n_0_1702;
   wire n_0_1703;
   wire n_0_1704;
   wire n_0_1705;
   wire n_0_1706;
   wire n_0_1707;
   wire n_0_1708;
   wire n_0_1709;
   wire n_0_1710;
   wire n_0_1711;
   wire n_0_1712;
   wire n_0_1713;
   wire n_0_1714;
   wire n_0_1715;
   wire n_0_1716;
   wire n_0_1717;
   wire n_0_1718;
   wire n_0_1719;
   wire n_0_1720;
   wire n_0_1721;
   wire n_0_1722;
   wire n_0_1723;
   wire n_0_1724;
   wire n_0_1725;
   wire n_0_1726;
   wire n_0_1727;
   wire n_0_1728;
   wire n_0_1729;
   wire n_0_1730;
   wire n_0_1731;
   wire n_0_1732;
   wire n_0_1733;
   wire n_0_1734;
   wire n_0_1735;
   wire n_0_1736;
   wire n_0_1737;
   wire n_0_1738;
   wire n_0_1739;
   wire n_0_1740;
   wire n_0_1741;
   wire n_0_1742;
   wire n_0_1743;
   wire n_0_1744;
   wire n_0_1745;
   wire n_0_1746;
   wire n_0_1747;
   wire n_0_1748;
   wire n_0_1749;
   wire n_0_1750;
   wire n_0_1751;
   wire n_0_1752;
   wire n_0_1753;
   wire n_0_1754;
   wire n_0_1755;
   wire n_0_1756;
   wire n_0_1757;
   wire n_0_1758;
   wire n_0_1759;
   wire n_0_1760;
   wire n_0_72_0;
   wire n_0_1762;
   wire n_0_1763;
   wire n_0_1761;
   wire n_0_73_0;
   wire n_0_73_1;
   wire n_0_1764;
   wire n_0_73_2;
   wire n_0_1765;
   wire n_0_73_3;
   wire n_0_1766;
   wire n_0_73_4;
   wire n_0_1767;
   wire n_0_73_5;
   wire n_0_1768;
   wire n_0_73_6;
   wire n_0_1769;
   wire n_0_73_7;
   wire n_0_1770;
   wire n_0_73_8;
   wire n_0_1771;
   wire n_0_73_9;
   wire n_0_1772;
   wire n_0_73_10;
   wire n_0_1773;
   wire n_0_73_11;
   wire n_0_1774;
   wire n_0_73_12;
   wire n_0_1775;
   wire n_0_73_13;
   wire n_0_1776;
   wire n_0_73_14;
   wire n_0_1777;
   wire n_0_73_15;
   wire n_0_1778;
   wire n_0_73_16;
   wire n_0_1779;
   wire n_0_73_17;
   wire n_0_1780;
   wire n_0_73_18;
   wire n_0_1781;
   wire n_0_73_19;
   wire n_0_1782;
   wire n_0_73_20;
   wire n_0_1783;
   wire n_0_73_21;
   wire n_0_1784;
   wire n_0_73_22;
   wire n_0_1785;
   wire n_0_73_23;
   wire n_0_1786;
   wire n_0_73_24;
   wire n_0_1787;
   wire n_0_73_25;
   wire n_0_1788;
   wire n_0_73_26;
   wire n_0_1789;
   wire n_0_73_27;
   wire n_0_1790;
   wire n_0_73_28;
   wire n_0_1791;
   wire n_0_73_29;
   wire n_0_1792;
   wire n_0_73_30;
   wire n_0_73_31;
   wire n_0_1793;
   wire n_0_73_32;
   wire n_0_1794;
   wire n_0_1795;
   wire n_0_1796;
   wire n_0_1797;
   wire n_0_1798;
   wire n_0_1799;
   wire n_0_1800;
   wire n_0_1801;
   wire n_0_1802;
   wire n_0_1803;
   wire n_0_1804;
   wire n_0_1805;
   wire n_0_1806;
   wire n_0_1807;
   wire n_0_1808;
   wire n_0_1809;
   wire n_0_1810;
   wire n_0_1811;
   wire n_0_1812;
   wire n_0_1813;
   wire n_0_1814;
   wire n_0_1815;
   wire n_0_1816;
   wire n_0_1817;
   wire n_0_1818;
   wire n_0_1819;
   wire n_0_1820;
   wire n_0_1821;
   wire n_0_1822;
   wire n_0_1823;
   wire n_0_1824;
   wire n_0_1825;
   wire n_0_1826;
   wire n_0_1827;
   wire n_0_1828;
   wire n_0_1829;
   wire n_0_1830;
   wire n_0_1831;
   wire n_0_1832;
   wire n_0_1833;
   wire n_0_1834;
   wire n_0_1835;
   wire n_0_1836;
   wire n_0_1837;
   wire n_0_1838;
   wire n_0_1839;
   wire n_0_1840;
   wire n_0_1841;
   wire n_0_1842;
   wire n_0_1843;
   wire n_0_1844;
   wire n_0_1845;
   wire n_0_1846;
   wire n_0_1847;
   wire n_0_1848;
   wire n_0_1849;
   wire n_0_1850;
   wire n_0_1851;
   wire n_0_1852;
   wire n_0_1853;
   wire n_0_1854;
   wire n_0_1855;
   wire n_0_1856;
   wire n_0_1857;
   wire n_0_1858;
   wire n_0_76_0;
   wire n_0_1860;
   wire n_0_1861;
   wire n_0_1859;
   wire n_0_77_0;
   wire n_0_77_1;
   wire n_0_1862;
   wire n_0_77_2;
   wire n_0_1863;
   wire n_0_77_3;
   wire n_0_1864;
   wire n_0_77_4;
   wire n_0_1865;
   wire n_0_77_5;
   wire n_0_1866;
   wire n_0_77_6;
   wire n_0_1867;
   wire n_0_77_7;
   wire n_0_1868;
   wire n_0_77_8;
   wire n_0_1869;
   wire n_0_77_9;
   wire n_0_1870;
   wire n_0_77_10;
   wire n_0_1871;
   wire n_0_77_11;
   wire n_0_1872;
   wire n_0_77_12;
   wire n_0_1873;
   wire n_0_77_13;
   wire n_0_1874;
   wire n_0_77_14;
   wire n_0_1875;
   wire n_0_77_15;
   wire n_0_1876;
   wire n_0_77_16;
   wire n_0_1877;
   wire n_0_77_17;
   wire n_0_1878;
   wire n_0_77_18;
   wire n_0_1879;
   wire n_0_77_19;
   wire n_0_1880;
   wire n_0_77_20;
   wire n_0_1881;
   wire n_0_77_21;
   wire n_0_1882;
   wire n_0_77_22;
   wire n_0_1883;
   wire n_0_77_23;
   wire n_0_1884;
   wire n_0_77_24;
   wire n_0_1885;
   wire n_0_77_25;
   wire n_0_1886;
   wire n_0_77_26;
   wire n_0_1887;
   wire n_0_77_27;
   wire n_0_1888;
   wire n_0_77_28;
   wire n_0_1889;
   wire n_0_77_29;
   wire n_0_1890;
   wire n_0_77_30;
   wire n_0_77_31;
   wire n_0_1891;
   wire n_0_77_32;
   wire n_0_1892;
   wire n_0_1893;
   wire n_0_1894;
   wire n_0_1895;
   wire n_0_1896;
   wire n_0_1897;
   wire n_0_1898;
   wire n_0_1899;
   wire n_0_1900;
   wire n_0_1901;
   wire n_0_1902;
   wire n_0_1903;
   wire n_0_1904;
   wire n_0_1905;
   wire n_0_1906;
   wire n_0_1907;
   wire n_0_1908;
   wire n_0_1909;
   wire n_0_1910;
   wire n_0_1911;
   wire n_0_1912;
   wire n_0_1913;
   wire n_0_1914;
   wire n_0_1915;
   wire n_0_1916;
   wire n_0_1917;
   wire n_0_1918;
   wire n_0_1919;
   wire n_0_1920;
   wire n_0_1921;
   wire n_0_1922;
   wire n_0_1923;
   wire n_0_1924;
   wire n_0_1925;
   wire n_0_1926;
   wire n_0_1927;
   wire n_0_1928;
   wire n_0_1929;
   wire n_0_1930;
   wire n_0_1931;
   wire n_0_1932;
   wire n_0_1933;
   wire n_0_1934;
   wire n_0_1935;
   wire n_0_1936;
   wire n_0_1937;
   wire n_0_1938;
   wire n_0_1939;
   wire n_0_1940;
   wire n_0_1941;
   wire n_0_1942;
   wire n_0_1943;
   wire n_0_1944;
   wire n_0_1945;
   wire n_0_1946;
   wire n_0_1947;
   wire n_0_1948;
   wire n_0_1949;
   wire n_0_1950;
   wire n_0_1951;
   wire n_0_1952;
   wire n_0_1953;
   wire n_0_1954;
   wire n_0_1955;
   wire n_0_1956;
   wire n_0_80_0;
   wire n_0_1958;
   wire n_0_1959;
   wire n_0_1957;
   wire n_0_81_0;
   wire n_0_81_1;
   wire n_0_1960;
   wire n_0_81_2;
   wire n_0_1961;
   wire n_0_81_3;
   wire n_0_1962;
   wire n_0_81_4;
   wire n_0_1963;
   wire n_0_81_5;
   wire n_0_1964;
   wire n_0_81_6;
   wire n_0_1965;
   wire n_0_81_7;
   wire n_0_1966;
   wire n_0_81_8;
   wire n_0_1967;
   wire n_0_81_9;
   wire n_0_1968;
   wire n_0_81_10;
   wire n_0_1969;
   wire n_0_81_11;
   wire n_0_1970;
   wire n_0_81_12;
   wire n_0_1971;
   wire n_0_81_13;
   wire n_0_1972;
   wire n_0_81_14;
   wire n_0_1973;
   wire n_0_81_15;
   wire n_0_1974;
   wire n_0_81_16;
   wire n_0_1975;
   wire n_0_81_17;
   wire n_0_1976;
   wire n_0_81_18;
   wire n_0_1977;
   wire n_0_81_19;
   wire n_0_1978;
   wire n_0_81_20;
   wire n_0_1979;
   wire n_0_81_21;
   wire n_0_1980;
   wire n_0_81_22;
   wire n_0_1981;
   wire n_0_81_23;
   wire n_0_1982;
   wire n_0_81_24;
   wire n_0_1983;
   wire n_0_81_25;
   wire n_0_1984;
   wire n_0_81_26;
   wire n_0_1985;
   wire n_0_81_27;
   wire n_0_1986;
   wire n_0_81_28;
   wire n_0_1987;
   wire n_0_81_29;
   wire n_0_1988;
   wire n_0_81_30;
   wire n_0_81_31;
   wire n_0_1989;
   wire n_0_81_32;
   wire n_0_1990;
   wire n_0_1991;
   wire n_0_1992;
   wire n_0_1993;
   wire n_0_1994;
   wire n_0_1995;
   wire n_0_1996;
   wire n_0_1997;
   wire n_0_1998;
   wire n_0_1999;
   wire n_0_2000;
   wire n_0_2001;
   wire n_0_2002;
   wire n_0_2003;
   wire n_0_2004;
   wire n_0_2005;
   wire n_0_2006;
   wire n_0_2007;
   wire n_0_2008;
   wire n_0_2009;
   wire n_0_2010;
   wire n_0_2011;
   wire n_0_2012;
   wire n_0_2013;
   wire n_0_2014;
   wire n_0_2015;
   wire n_0_2016;
   wire n_0_2017;
   wire n_0_2018;
   wire n_0_2019;
   wire n_0_2020;
   wire n_0_2021;
   wire n_0_2022;
   wire n_0_2023;
   wire n_0_2024;
   wire n_0_2025;
   wire n_0_2026;
   wire n_0_2027;
   wire n_0_2028;
   wire n_0_2029;
   wire n_0_2030;
   wire n_0_2031;
   wire n_0_2032;
   wire n_0_2033;
   wire n_0_2034;
   wire n_0_2035;
   wire n_0_2036;
   wire n_0_2037;
   wire n_0_2038;
   wire n_0_2039;
   wire n_0_2040;
   wire n_0_2041;
   wire n_0_2042;
   wire n_0_2043;
   wire n_0_2044;
   wire n_0_2045;
   wire n_0_2046;
   wire n_0_2047;
   wire n_0_2048;
   wire n_0_2049;
   wire n_0_2050;
   wire n_0_2051;
   wire n_0_2052;
   wire n_0_2053;
   wire n_0_2054;
   wire n_0_84_0;
   wire n_0_2056;
   wire n_0_2057;
   wire n_0_2055;
   wire n_0_85_0;
   wire n_0_85_1;
   wire n_0_2058;
   wire n_0_85_2;
   wire n_0_2059;
   wire n_0_85_3;
   wire n_0_2060;
   wire n_0_85_4;
   wire n_0_2061;
   wire n_0_85_5;
   wire n_0_2062;
   wire n_0_85_6;
   wire n_0_2063;
   wire n_0_85_7;
   wire n_0_2064;
   wire n_0_85_8;
   wire n_0_2065;
   wire n_0_85_9;
   wire n_0_2066;
   wire n_0_85_10;
   wire n_0_2067;
   wire n_0_85_11;
   wire n_0_2068;
   wire n_0_85_12;
   wire n_0_2069;
   wire n_0_85_13;
   wire n_0_2070;
   wire n_0_85_14;
   wire n_0_2071;
   wire n_0_85_15;
   wire n_0_2072;
   wire n_0_85_16;
   wire n_0_2073;
   wire n_0_85_17;
   wire n_0_2074;
   wire n_0_85_18;
   wire n_0_2075;
   wire n_0_85_19;
   wire n_0_2076;
   wire n_0_85_20;
   wire n_0_2077;
   wire n_0_85_21;
   wire n_0_2078;
   wire n_0_85_22;
   wire n_0_2079;
   wire n_0_85_23;
   wire n_0_2080;
   wire n_0_85_24;
   wire n_0_2081;
   wire n_0_85_25;
   wire n_0_2082;
   wire n_0_85_26;
   wire n_0_2083;
   wire n_0_85_27;
   wire n_0_2084;
   wire n_0_85_28;
   wire n_0_2085;
   wire n_0_85_29;
   wire n_0_2086;
   wire n_0_85_30;
   wire n_0_85_31;
   wire n_0_2087;
   wire n_0_85_32;
   wire n_0_2088;
   wire n_0_2089;
   wire n_0_2090;
   wire n_0_2091;
   wire n_0_2092;
   wire n_0_2093;
   wire n_0_2094;
   wire n_0_2095;
   wire n_0_2096;
   wire n_0_2097;
   wire n_0_2098;
   wire n_0_2099;
   wire n_0_2100;
   wire n_0_2101;
   wire n_0_2102;
   wire n_0_2103;
   wire n_0_2104;
   wire n_0_2105;
   wire n_0_2106;
   wire n_0_2107;
   wire n_0_2108;
   wire n_0_2109;
   wire n_0_2110;
   wire n_0_2111;
   wire n_0_2112;
   wire n_0_2113;
   wire n_0_2114;
   wire n_0_2115;
   wire n_0_2116;
   wire n_0_2117;
   wire n_0_2118;
   wire n_0_2119;
   wire n_0_2120;
   wire n_0_2121;
   wire n_0_2122;
   wire n_0_2123;
   wire n_0_2124;
   wire n_0_2125;
   wire n_0_2126;
   wire n_0_2127;
   wire n_0_2128;
   wire n_0_2129;
   wire n_0_2130;
   wire n_0_2131;
   wire n_0_2132;
   wire n_0_2133;
   wire n_0_2134;
   wire n_0_2135;
   wire n_0_2136;
   wire n_0_2137;
   wire n_0_2138;
   wire n_0_2139;
   wire n_0_2140;
   wire n_0_2141;
   wire n_0_2142;
   wire n_0_2143;
   wire n_0_2144;
   wire n_0_2145;
   wire n_0_2146;
   wire n_0_2147;
   wire n_0_2148;
   wire n_0_2149;
   wire n_0_2150;
   wire n_0_2151;
   wire n_0_2152;
   wire n_0_88_0;
   wire n_0_2154;
   wire n_0_2155;
   wire n_0_2153;
   wire n_0_89_0;
   wire n_0_89_1;
   wire n_0_2156;
   wire n_0_89_2;
   wire n_0_2157;
   wire n_0_89_3;
   wire n_0_2158;
   wire n_0_89_4;
   wire n_0_2159;
   wire n_0_89_5;
   wire n_0_2160;
   wire n_0_89_6;
   wire n_0_2161;
   wire n_0_89_7;
   wire n_0_2162;
   wire n_0_89_8;
   wire n_0_2163;
   wire n_0_89_9;
   wire n_0_2164;
   wire n_0_89_10;
   wire n_0_2165;
   wire n_0_89_11;
   wire n_0_2166;
   wire n_0_89_12;
   wire n_0_2167;
   wire n_0_89_13;
   wire n_0_2168;
   wire n_0_89_14;
   wire n_0_2169;
   wire n_0_89_15;
   wire n_0_2170;
   wire n_0_89_16;
   wire n_0_2171;
   wire n_0_89_17;
   wire n_0_2172;
   wire n_0_89_18;
   wire n_0_2173;
   wire n_0_89_19;
   wire n_0_2174;
   wire n_0_89_20;
   wire n_0_2175;
   wire n_0_89_21;
   wire n_0_2176;
   wire n_0_89_22;
   wire n_0_2177;
   wire n_0_89_23;
   wire n_0_2178;
   wire n_0_89_24;
   wire n_0_2179;
   wire n_0_89_25;
   wire n_0_2180;
   wire n_0_89_26;
   wire n_0_2181;
   wire n_0_89_27;
   wire n_0_2182;
   wire n_0_89_28;
   wire n_0_2183;
   wire n_0_89_29;
   wire n_0_2184;
   wire n_0_89_30;
   wire n_0_89_31;
   wire n_0_2185;
   wire n_0_89_32;
   wire n_0_2186;
   wire n_0_2187;
   wire n_0_2188;
   wire n_0_2189;
   wire n_0_2190;
   wire n_0_2191;
   wire n_0_2192;
   wire n_0_2193;
   wire n_0_2194;
   wire n_0_2195;
   wire n_0_2196;
   wire n_0_2197;
   wire n_0_2198;
   wire n_0_2199;
   wire n_0_2200;
   wire n_0_2201;
   wire n_0_2202;
   wire n_0_2203;
   wire n_0_2204;
   wire n_0_2205;
   wire n_0_2206;
   wire n_0_2207;
   wire n_0_2208;
   wire n_0_2209;
   wire n_0_2210;
   wire n_0_2211;
   wire n_0_2212;
   wire n_0_2213;
   wire n_0_2214;
   wire n_0_2215;
   wire n_0_2216;
   wire n_0_2217;
   wire n_0_2218;
   wire n_0_2219;
   wire n_0_2220;
   wire n_0_2221;
   wire n_0_2222;
   wire n_0_2223;
   wire n_0_2224;
   wire n_0_2225;
   wire n_0_2226;
   wire n_0_2227;
   wire n_0_2228;
   wire n_0_2229;
   wire n_0_2230;
   wire n_0_2231;
   wire n_0_2232;
   wire n_0_2233;
   wire n_0_2234;
   wire n_0_2235;
   wire n_0_2236;
   wire n_0_2237;
   wire n_0_2238;
   wire n_0_2239;
   wire n_0_2240;
   wire n_0_2241;
   wire n_0_2242;
   wire n_0_2243;
   wire n_0_2244;
   wire n_0_2245;
   wire n_0_2246;
   wire n_0_2247;
   wire n_0_2248;
   wire n_0_2249;
   wire n_0_2250;
   wire n_0_92_0;
   wire n_0_2252;
   wire n_0_2253;
   wire n_0_2251;
   wire n_0_93_0;
   wire n_0_93_1;
   wire n_0_2254;
   wire n_0_93_2;
   wire n_0_2255;
   wire n_0_93_3;
   wire n_0_2256;
   wire n_0_93_4;
   wire n_0_2257;
   wire n_0_93_5;
   wire n_0_2258;
   wire n_0_93_6;
   wire n_0_2259;
   wire n_0_93_7;
   wire n_0_2260;
   wire n_0_93_8;
   wire n_0_2261;
   wire n_0_93_9;
   wire n_0_2262;
   wire n_0_93_10;
   wire n_0_2263;
   wire n_0_93_11;
   wire n_0_2264;
   wire n_0_93_12;
   wire n_0_2265;
   wire n_0_93_13;
   wire n_0_2266;
   wire n_0_93_14;
   wire n_0_2267;
   wire n_0_93_15;
   wire n_0_2268;
   wire n_0_93_16;
   wire n_0_2269;
   wire n_0_93_17;
   wire n_0_2270;
   wire n_0_93_18;
   wire n_0_2271;
   wire n_0_93_19;
   wire n_0_2272;
   wire n_0_93_20;
   wire n_0_2273;
   wire n_0_93_21;
   wire n_0_2274;
   wire n_0_93_22;
   wire n_0_2275;
   wire n_0_93_23;
   wire n_0_2276;
   wire n_0_93_24;
   wire n_0_2277;
   wire n_0_93_25;
   wire n_0_2278;
   wire n_0_93_26;
   wire n_0_2279;
   wire n_0_93_27;
   wire n_0_2280;
   wire n_0_93_28;
   wire n_0_2281;
   wire n_0_93_29;
   wire n_0_2282;
   wire n_0_93_30;
   wire n_0_93_31;
   wire n_0_2283;
   wire n_0_93_32;
   wire n_0_2284;
   wire n_0_2285;
   wire n_0_2286;
   wire n_0_2287;
   wire n_0_2288;
   wire n_0_2289;
   wire n_0_2290;
   wire n_0_2291;
   wire n_0_2292;
   wire n_0_2293;
   wire n_0_2294;
   wire n_0_2295;
   wire n_0_2296;
   wire n_0_2297;
   wire n_0_2298;
   wire n_0_2299;
   wire n_0_2300;
   wire n_0_2301;
   wire n_0_2302;
   wire n_0_2303;
   wire n_0_2304;
   wire n_0_2305;
   wire n_0_2306;
   wire n_0_2307;
   wire n_0_2308;
   wire n_0_2309;
   wire n_0_2310;
   wire n_0_2311;
   wire n_0_2312;
   wire n_0_2313;
   wire n_0_2314;
   wire n_0_2315;
   wire n_0_2316;
   wire n_0_2317;
   wire n_0_2318;
   wire n_0_2319;
   wire n_0_2320;
   wire n_0_2321;
   wire n_0_2322;
   wire n_0_2323;
   wire n_0_2324;
   wire n_0_2325;
   wire n_0_2326;
   wire n_0_2327;
   wire n_0_2328;
   wire n_0_2329;
   wire n_0_2330;
   wire n_0_2331;
   wire n_0_2332;
   wire n_0_2333;
   wire n_0_2334;
   wire n_0_2335;
   wire n_0_2336;
   wire n_0_2337;
   wire n_0_2338;
   wire n_0_2339;
   wire n_0_2340;
   wire n_0_2341;
   wire n_0_2342;
   wire n_0_2343;
   wire n_0_2344;
   wire n_0_2345;
   wire n_0_2346;
   wire n_0_2347;
   wire n_0_2348;
   wire n_0_96_0;
   wire n_0_2350;
   wire n_0_2351;
   wire n_0_2349;
   wire n_0_97_0;
   wire n_0_97_1;
   wire n_0_2352;
   wire n_0_97_2;
   wire n_0_2353;
   wire n_0_97_3;
   wire n_0_2354;
   wire n_0_97_4;
   wire n_0_2355;
   wire n_0_97_5;
   wire n_0_2356;
   wire n_0_97_6;
   wire n_0_2357;
   wire n_0_97_7;
   wire n_0_2358;
   wire n_0_97_8;
   wire n_0_2359;
   wire n_0_97_9;
   wire n_0_2360;
   wire n_0_97_10;
   wire n_0_2361;
   wire n_0_97_11;
   wire n_0_2362;
   wire n_0_97_12;
   wire n_0_2363;
   wire n_0_97_13;
   wire n_0_2364;
   wire n_0_97_14;
   wire n_0_2365;
   wire n_0_97_15;
   wire n_0_2366;
   wire n_0_97_16;
   wire n_0_2367;
   wire n_0_97_17;
   wire n_0_2368;
   wire n_0_97_18;
   wire n_0_2369;
   wire n_0_97_19;
   wire n_0_2370;
   wire n_0_97_20;
   wire n_0_2371;
   wire n_0_97_21;
   wire n_0_2372;
   wire n_0_97_22;
   wire n_0_2373;
   wire n_0_97_23;
   wire n_0_2374;
   wire n_0_97_24;
   wire n_0_2375;
   wire n_0_97_25;
   wire n_0_2376;
   wire n_0_97_26;
   wire n_0_2377;
   wire n_0_97_27;
   wire n_0_2378;
   wire n_0_97_28;
   wire n_0_2379;
   wire n_0_97_29;
   wire n_0_2380;
   wire n_0_97_30;
   wire n_0_97_31;
   wire n_0_2381;
   wire n_0_97_32;
   wire n_0_2382;
   wire n_0_2383;
   wire n_0_2384;
   wire n_0_2385;
   wire n_0_2386;
   wire n_0_2387;
   wire n_0_2388;
   wire n_0_2389;
   wire n_0_2390;
   wire n_0_2391;
   wire n_0_2392;
   wire n_0_2393;
   wire n_0_2394;
   wire n_0_2395;
   wire n_0_2396;
   wire n_0_2397;
   wire n_0_2398;
   wire n_0_2399;
   wire n_0_2400;
   wire n_0_2401;
   wire n_0_2402;
   wire n_0_2403;
   wire n_0_2404;
   wire n_0_2405;
   wire n_0_2406;
   wire n_0_2407;
   wire n_0_2408;
   wire n_0_2409;
   wire n_0_2410;
   wire n_0_2411;
   wire n_0_2412;
   wire n_0_2413;
   wire n_0_2414;
   wire n_0_2415;
   wire n_0_2416;
   wire n_0_2417;
   wire n_0_2418;
   wire n_0_2419;
   wire n_0_2420;
   wire n_0_2421;
   wire n_0_2422;
   wire n_0_2423;
   wire n_0_2424;
   wire n_0_2425;
   wire n_0_2426;
   wire n_0_2427;
   wire n_0_2428;
   wire n_0_2429;
   wire n_0_2430;
   wire n_0_2431;
   wire n_0_2432;
   wire n_0_2433;
   wire n_0_2434;
   wire n_0_2435;
   wire n_0_2436;
   wire n_0_2437;
   wire n_0_2438;
   wire n_0_2439;
   wire n_0_2440;
   wire n_0_2441;
   wire n_0_2442;
   wire n_0_2443;
   wire n_0_2444;
   wire n_0_2445;
   wire n_0_2446;
   wire n_0_100_0;
   wire n_0_2448;
   wire n_0_2449;
   wire n_0_2447;
   wire n_0_101_0;
   wire n_0_101_1;
   wire n_0_2450;
   wire n_0_101_2;
   wire n_0_2451;
   wire n_0_101_3;
   wire n_0_2452;
   wire n_0_101_4;
   wire n_0_2453;
   wire n_0_101_5;
   wire n_0_2454;
   wire n_0_101_6;
   wire n_0_2455;
   wire n_0_101_7;
   wire n_0_2456;
   wire n_0_101_8;
   wire n_0_2457;
   wire n_0_101_9;
   wire n_0_2458;
   wire n_0_101_10;
   wire n_0_2459;
   wire n_0_101_11;
   wire n_0_2460;
   wire n_0_101_12;
   wire n_0_2461;
   wire n_0_101_13;
   wire n_0_2462;
   wire n_0_101_14;
   wire n_0_2463;
   wire n_0_101_15;
   wire n_0_2464;
   wire n_0_101_16;
   wire n_0_2465;
   wire n_0_101_17;
   wire n_0_2466;
   wire n_0_101_18;
   wire n_0_2467;
   wire n_0_101_19;
   wire n_0_2468;
   wire n_0_101_20;
   wire n_0_2469;
   wire n_0_101_21;
   wire n_0_2470;
   wire n_0_101_22;
   wire n_0_2471;
   wire n_0_101_23;
   wire n_0_2472;
   wire n_0_101_24;
   wire n_0_2473;
   wire n_0_101_25;
   wire n_0_2474;
   wire n_0_101_26;
   wire n_0_2475;
   wire n_0_101_27;
   wire n_0_2476;
   wire n_0_101_28;
   wire n_0_2477;
   wire n_0_101_29;
   wire n_0_2478;
   wire n_0_101_30;
   wire n_0_101_31;
   wire n_0_2479;
   wire n_0_101_32;
   wire n_0_2480;
   wire n_0_2481;
   wire n_0_2482;
   wire n_0_2483;
   wire n_0_2484;
   wire n_0_2485;
   wire n_0_2486;
   wire n_0_2487;
   wire n_0_2488;
   wire n_0_2489;
   wire n_0_2490;
   wire n_0_2491;
   wire n_0_2492;
   wire n_0_2493;
   wire n_0_2494;
   wire n_0_2495;
   wire n_0_2496;
   wire n_0_2497;
   wire n_0_2498;
   wire n_0_2499;
   wire n_0_2500;
   wire n_0_2501;
   wire n_0_2502;
   wire n_0_2503;
   wire n_0_2504;
   wire n_0_2505;
   wire n_0_2506;
   wire n_0_2507;
   wire n_0_2508;
   wire n_0_2509;
   wire n_0_2510;
   wire n_0_2511;
   wire n_0_2512;
   wire n_0_2513;
   wire n_0_2514;
   wire n_0_2515;
   wire n_0_2516;
   wire n_0_2517;
   wire n_0_2518;
   wire n_0_2519;
   wire n_0_2520;
   wire n_0_2521;
   wire n_0_2522;
   wire n_0_2523;
   wire n_0_2524;
   wire n_0_2525;
   wire n_0_2526;
   wire n_0_2527;
   wire n_0_2528;
   wire n_0_2529;
   wire n_0_2530;
   wire n_0_2531;
   wire n_0_2532;
   wire n_0_2533;
   wire n_0_2534;
   wire n_0_2535;
   wire n_0_2536;
   wire n_0_2537;
   wire n_0_2538;
   wire n_0_2539;
   wire n_0_2540;
   wire n_0_2541;
   wire n_0_2542;
   wire n_0_2543;
   wire n_0_2544;
   wire n_0_104_0;
   wire n_0_2546;
   wire n_0_2547;
   wire n_0_2545;
   wire n_0_105_0;
   wire n_0_105_1;
   wire n_0_2548;
   wire n_0_105_2;
   wire n_0_2549;
   wire n_0_105_3;
   wire n_0_2550;
   wire n_0_105_4;
   wire n_0_2551;
   wire n_0_105_5;
   wire n_0_2552;
   wire n_0_105_6;
   wire n_0_2553;
   wire n_0_105_7;
   wire n_0_2554;
   wire n_0_105_8;
   wire n_0_2555;
   wire n_0_105_9;
   wire n_0_2556;
   wire n_0_105_10;
   wire n_0_2557;
   wire n_0_105_11;
   wire n_0_2558;
   wire n_0_105_12;
   wire n_0_2559;
   wire n_0_105_13;
   wire n_0_2560;
   wire n_0_105_14;
   wire n_0_2561;
   wire n_0_105_15;
   wire n_0_2562;
   wire n_0_105_16;
   wire n_0_2563;
   wire n_0_105_17;
   wire n_0_2564;
   wire n_0_105_18;
   wire n_0_2565;
   wire n_0_105_19;
   wire n_0_2566;
   wire n_0_105_20;
   wire n_0_2567;
   wire n_0_105_21;
   wire n_0_2568;
   wire n_0_105_22;
   wire n_0_2569;
   wire n_0_105_23;
   wire n_0_2570;
   wire n_0_105_24;
   wire n_0_2571;
   wire n_0_105_25;
   wire n_0_2572;
   wire n_0_105_26;
   wire n_0_2573;
   wire n_0_105_27;
   wire n_0_2574;
   wire n_0_105_28;
   wire n_0_2575;
   wire n_0_105_29;
   wire n_0_2576;
   wire n_0_105_30;
   wire n_0_105_31;
   wire n_0_2577;
   wire n_0_105_32;
   wire n_0_2578;
   wire n_0_2579;
   wire n_0_2580;
   wire n_0_2581;
   wire n_0_2582;
   wire n_0_2583;
   wire n_0_2584;
   wire n_0_2585;
   wire n_0_2586;
   wire n_0_2587;
   wire n_0_2588;
   wire n_0_2589;
   wire n_0_2590;
   wire n_0_2591;
   wire n_0_2592;
   wire n_0_2593;
   wire n_0_2594;
   wire n_0_2595;
   wire n_0_2596;
   wire n_0_2597;
   wire n_0_2598;
   wire n_0_2599;
   wire n_0_2600;
   wire n_0_2601;
   wire n_0_2602;
   wire n_0_2603;
   wire n_0_2604;
   wire n_0_2605;
   wire n_0_2606;
   wire n_0_2607;
   wire n_0_2608;
   wire n_0_2609;
   wire n_0_2610;
   wire n_0_2611;
   wire n_0_2612;
   wire n_0_2613;
   wire n_0_2614;
   wire n_0_2615;
   wire n_0_2616;
   wire n_0_2617;
   wire n_0_2618;
   wire n_0_2619;
   wire n_0_2620;
   wire n_0_2621;
   wire n_0_2622;
   wire n_0_2623;
   wire n_0_2624;
   wire n_0_2625;
   wire n_0_2626;
   wire n_0_2627;
   wire n_0_2628;
   wire n_0_2629;
   wire n_0_2630;
   wire n_0_2631;
   wire n_0_2632;
   wire n_0_2633;
   wire n_0_2634;
   wire n_0_2635;
   wire n_0_2636;
   wire n_0_2637;
   wire n_0_2638;
   wire n_0_2639;
   wire n_0_2640;
   wire n_0_2641;
   wire n_0_2642;
   wire n_0_108_0;
   wire n_0_2644;
   wire n_0_2645;
   wire n_0_2643;
   wire n_0_109_0;
   wire n_0_109_1;
   wire n_0_2646;
   wire n_0_109_2;
   wire n_0_2647;
   wire n_0_109_3;
   wire n_0_2648;
   wire n_0_109_4;
   wire n_0_2649;
   wire n_0_109_5;
   wire n_0_2650;
   wire n_0_109_6;
   wire n_0_2651;
   wire n_0_109_7;
   wire n_0_2652;
   wire n_0_109_8;
   wire n_0_2653;
   wire n_0_109_9;
   wire n_0_2654;
   wire n_0_109_10;
   wire n_0_2655;
   wire n_0_109_11;
   wire n_0_2656;
   wire n_0_109_12;
   wire n_0_2657;
   wire n_0_109_13;
   wire n_0_2658;
   wire n_0_109_14;
   wire n_0_2659;
   wire n_0_109_15;
   wire n_0_2660;
   wire n_0_109_16;
   wire n_0_2661;
   wire n_0_109_17;
   wire n_0_2662;
   wire n_0_109_18;
   wire n_0_2663;
   wire n_0_109_19;
   wire n_0_2664;
   wire n_0_109_20;
   wire n_0_2665;
   wire n_0_109_21;
   wire n_0_2666;
   wire n_0_109_22;
   wire n_0_2667;
   wire n_0_109_23;
   wire n_0_2668;
   wire n_0_109_24;
   wire n_0_2669;
   wire n_0_109_25;
   wire n_0_2670;
   wire n_0_109_26;
   wire n_0_2671;
   wire n_0_109_27;
   wire n_0_2672;
   wire n_0_109_28;
   wire n_0_2673;
   wire n_0_109_29;
   wire n_0_2674;
   wire n_0_109_30;
   wire n_0_109_31;
   wire n_0_2675;
   wire n_0_109_32;
   wire n_0_2676;
   wire n_0_2677;
   wire n_0_2678;
   wire n_0_2679;
   wire n_0_2680;
   wire n_0_2681;
   wire n_0_2682;
   wire n_0_2683;
   wire n_0_2684;
   wire n_0_2685;
   wire n_0_2686;
   wire n_0_2687;
   wire n_0_2688;
   wire n_0_2689;
   wire n_0_2690;
   wire n_0_2691;
   wire n_0_2692;
   wire n_0_2693;
   wire n_0_2694;
   wire n_0_2695;
   wire n_0_2696;
   wire n_0_2697;
   wire n_0_2698;
   wire n_0_2699;
   wire n_0_2700;
   wire n_0_2701;
   wire n_0_2702;
   wire n_0_2703;
   wire n_0_2704;
   wire n_0_2705;
   wire n_0_2706;
   wire n_0_2707;
   wire n_0_2708;
   wire n_0_2709;
   wire n_0_2710;
   wire n_0_2711;
   wire n_0_2712;
   wire n_0_2713;
   wire n_0_2714;
   wire n_0_2715;
   wire n_0_2716;
   wire n_0_2717;
   wire n_0_2718;
   wire n_0_2719;
   wire n_0_2720;
   wire n_0_2721;
   wire n_0_2722;
   wire n_0_2723;
   wire n_0_2724;
   wire n_0_2725;
   wire n_0_2726;
   wire n_0_2727;
   wire n_0_2728;
   wire n_0_2729;
   wire n_0_2730;
   wire n_0_2731;
   wire n_0_2732;
   wire n_0_2733;
   wire n_0_2734;
   wire n_0_2735;
   wire n_0_2736;
   wire n_0_2737;
   wire n_0_2738;
   wire n_0_2739;
   wire n_0_2740;
   wire n_0_112_0;
   wire n_0_2742;
   wire n_0_2743;
   wire n_0_2741;
   wire n_0_113_0;
   wire n_0_113_1;
   wire n_0_2744;
   wire n_0_113_2;
   wire n_0_2745;
   wire n_0_113_3;
   wire n_0_2746;
   wire n_0_113_4;
   wire n_0_2747;
   wire n_0_113_5;
   wire n_0_2748;
   wire n_0_113_6;
   wire n_0_2749;
   wire n_0_113_7;
   wire n_0_2750;
   wire n_0_113_8;
   wire n_0_2751;
   wire n_0_113_9;
   wire n_0_2752;
   wire n_0_113_10;
   wire n_0_2753;
   wire n_0_113_11;
   wire n_0_2754;
   wire n_0_113_12;
   wire n_0_2755;
   wire n_0_113_13;
   wire n_0_2756;
   wire n_0_113_14;
   wire n_0_2757;
   wire n_0_113_15;
   wire n_0_2758;
   wire n_0_113_16;
   wire n_0_2759;
   wire n_0_113_17;
   wire n_0_2760;
   wire n_0_113_18;
   wire n_0_2761;
   wire n_0_113_19;
   wire n_0_2762;
   wire n_0_113_20;
   wire n_0_2763;
   wire n_0_113_21;
   wire n_0_2764;
   wire n_0_113_22;
   wire n_0_2765;
   wire n_0_113_23;
   wire n_0_2766;
   wire n_0_113_24;
   wire n_0_2767;
   wire n_0_113_25;
   wire n_0_2768;
   wire n_0_113_26;
   wire n_0_2769;
   wire n_0_113_27;
   wire n_0_2770;
   wire n_0_113_28;
   wire n_0_2771;
   wire n_0_113_29;
   wire n_0_2772;
   wire n_0_113_30;
   wire n_0_113_31;
   wire n_0_2773;
   wire n_0_113_32;
   wire n_0_2774;
   wire n_0_2775;
   wire n_0_2776;
   wire n_0_2777;
   wire n_0_2778;
   wire n_0_2779;
   wire n_0_2780;
   wire n_0_2781;
   wire n_0_2782;
   wire n_0_2783;
   wire n_0_2784;
   wire n_0_2785;
   wire n_0_2786;
   wire n_0_2787;
   wire n_0_2788;
   wire n_0_2789;
   wire n_0_2790;
   wire n_0_2791;
   wire n_0_2792;
   wire n_0_2793;
   wire n_0_2794;
   wire n_0_2795;
   wire n_0_2796;
   wire n_0_2797;
   wire n_0_2798;
   wire n_0_2799;
   wire n_0_2800;
   wire n_0_2801;
   wire n_0_2802;
   wire n_0_2803;
   wire n_0_2804;
   wire n_0_2805;
   wire n_0_2806;
   wire n_0_2807;
   wire n_0_2808;
   wire n_0_2809;
   wire n_0_2810;
   wire n_0_2811;
   wire n_0_2812;
   wire n_0_2813;
   wire n_0_2814;
   wire n_0_2815;
   wire n_0_2816;
   wire n_0_2817;
   wire n_0_2818;
   wire n_0_2819;
   wire n_0_2820;
   wire n_0_2821;
   wire n_0_2822;
   wire n_0_2823;
   wire n_0_2824;
   wire n_0_2825;
   wire n_0_2826;
   wire n_0_2827;
   wire n_0_2828;
   wire n_0_2829;
   wire n_0_2830;
   wire n_0_2831;
   wire n_0_2832;
   wire n_0_2833;
   wire n_0_2834;
   wire n_0_2835;
   wire n_0_2836;
   wire n_0_2837;
   wire n_0_2838;
   wire n_0_116_0;
   wire n_0_2840;
   wire n_0_2841;
   wire n_0_2839;
   wire n_0_117_0;
   wire n_0_117_1;
   wire n_0_2842;
   wire n_0_117_2;
   wire n_0_2843;
   wire n_0_117_3;
   wire n_0_2844;
   wire n_0_117_4;
   wire n_0_2845;
   wire n_0_117_5;
   wire n_0_2846;
   wire n_0_117_6;
   wire n_0_2847;
   wire n_0_117_7;
   wire n_0_2848;
   wire n_0_117_8;
   wire n_0_2849;
   wire n_0_117_9;
   wire n_0_2850;
   wire n_0_117_10;
   wire n_0_2851;
   wire n_0_117_11;
   wire n_0_2852;
   wire n_0_117_12;
   wire n_0_2853;
   wire n_0_117_13;
   wire n_0_2854;
   wire n_0_117_14;
   wire n_0_2855;
   wire n_0_117_15;
   wire n_0_2856;
   wire n_0_117_16;
   wire n_0_2857;
   wire n_0_117_17;
   wire n_0_2858;
   wire n_0_117_18;
   wire n_0_2859;
   wire n_0_117_19;
   wire n_0_2860;
   wire n_0_117_20;
   wire n_0_2861;
   wire n_0_117_21;
   wire n_0_2862;
   wire n_0_117_22;
   wire n_0_2863;
   wire n_0_117_23;
   wire n_0_2864;
   wire n_0_117_24;
   wire n_0_2865;
   wire n_0_117_25;
   wire n_0_2866;
   wire n_0_117_26;
   wire n_0_2867;
   wire n_0_117_27;
   wire n_0_2868;
   wire n_0_117_28;
   wire n_0_2869;
   wire n_0_117_29;
   wire n_0_2870;
   wire n_0_117_30;
   wire n_0_117_31;
   wire n_0_2871;
   wire n_0_117_32;
   wire n_0_2872;
   wire n_0_2873;
   wire n_0_2874;
   wire n_0_2875;
   wire n_0_2876;
   wire n_0_2877;
   wire n_0_2878;
   wire n_0_2879;
   wire n_0_2880;
   wire n_0_2881;
   wire n_0_2882;
   wire n_0_2883;
   wire n_0_2884;
   wire n_0_2885;
   wire n_0_2886;
   wire n_0_2887;
   wire n_0_2888;
   wire n_0_2889;
   wire n_0_2890;
   wire n_0_2891;
   wire n_0_2892;
   wire n_0_2893;
   wire n_0_2894;
   wire n_0_2895;
   wire n_0_2896;
   wire n_0_2897;
   wire n_0_2898;
   wire n_0_2899;
   wire n_0_2900;
   wire n_0_2901;
   wire n_0_2902;
   wire n_0_2903;
   wire n_0_2904;
   wire n_0_2905;
   wire n_0_2906;
   wire n_0_2907;
   wire n_0_2908;
   wire n_0_2909;
   wire n_0_2910;
   wire n_0_2911;
   wire n_0_2912;
   wire n_0_2913;
   wire n_0_2914;
   wire n_0_2915;
   wire n_0_2916;
   wire n_0_2917;
   wire n_0_2918;
   wire n_0_2919;
   wire n_0_2920;
   wire n_0_2921;
   wire n_0_2922;
   wire n_0_2923;
   wire n_0_2924;
   wire n_0_2925;
   wire n_0_2926;
   wire n_0_2927;
   wire n_0_2928;
   wire n_0_2929;
   wire n_0_2930;
   wire n_0_2931;
   wire n_0_2932;
   wire n_0_2933;
   wire n_0_2934;
   wire n_0_2935;
   wire n_0_2936;
   wire n_0_120_0;
   wire n_0_2938;
   wire n_0_2939;
   wire n_0_2937;
   wire n_0_121_0;
   wire n_0_121_1;
   wire n_0_2940;
   wire n_0_121_2;
   wire n_0_2941;
   wire n_0_121_3;
   wire n_0_2942;
   wire n_0_121_4;
   wire n_0_2943;
   wire n_0_121_5;
   wire n_0_2944;
   wire n_0_121_6;
   wire n_0_2945;
   wire n_0_121_7;
   wire n_0_2946;
   wire n_0_121_8;
   wire n_0_2947;
   wire n_0_121_9;
   wire n_0_2948;
   wire n_0_121_10;
   wire n_0_2949;
   wire n_0_121_11;
   wire n_0_2950;
   wire n_0_121_12;
   wire n_0_2951;
   wire n_0_121_13;
   wire n_0_2952;
   wire n_0_121_14;
   wire n_0_2953;
   wire n_0_121_15;
   wire n_0_2954;
   wire n_0_121_16;
   wire n_0_2955;
   wire n_0_121_17;
   wire n_0_2956;
   wire n_0_121_18;
   wire n_0_2957;
   wire n_0_121_19;
   wire n_0_2958;
   wire n_0_121_20;
   wire n_0_2959;
   wire n_0_121_21;
   wire n_0_2960;
   wire n_0_121_22;
   wire n_0_2961;
   wire n_0_121_23;
   wire n_0_2962;
   wire n_0_121_24;
   wire n_0_2963;
   wire n_0_121_25;
   wire n_0_2964;
   wire n_0_121_26;
   wire n_0_2965;
   wire n_0_121_27;
   wire n_0_2966;
   wire n_0_121_28;
   wire n_0_2967;
   wire n_0_121_29;
   wire n_0_2968;
   wire n_0_121_30;
   wire n_0_121_31;
   wire n_0_2969;
   wire n_0_121_32;
   wire n_0_2970;
   wire n_0_2971;
   wire n_0_2972;
   wire n_0_2973;
   wire n_0_2974;
   wire n_0_2975;
   wire n_0_2976;
   wire n_0_2977;
   wire n_0_2978;
   wire n_0_2979;
   wire n_0_2980;
   wire n_0_2981;
   wire n_0_2982;
   wire n_0_2983;
   wire n_0_2984;
   wire n_0_2985;
   wire n_0_2986;
   wire n_0_2987;
   wire n_0_2988;
   wire n_0_2989;
   wire n_0_2990;
   wire n_0_2991;
   wire n_0_2992;
   wire n_0_2993;
   wire n_0_2994;
   wire n_0_2995;
   wire n_0_2996;
   wire n_0_2997;
   wire n_0_2998;
   wire n_0_2999;
   wire n_0_3000;
   wire n_0_3001;
   wire n_0_3002;
   wire n_0_3003;
   wire n_0_3004;
   wire n_0_3005;
   wire n_0_3006;
   wire n_0_3007;
   wire n_0_3008;
   wire n_0_3009;
   wire n_0_3010;
   wire n_0_3011;
   wire n_0_3012;
   wire n_0_3013;
   wire n_0_3014;
   wire n_0_3015;
   wire n_0_3016;
   wire n_0_3017;
   wire n_0_3018;
   wire n_0_3019;
   wire n_0_3020;
   wire n_0_3021;
   wire n_0_3022;
   wire n_0_3023;
   wire n_0_3024;
   wire n_0_3025;
   wire n_0_3026;
   wire n_0_3027;
   wire n_0_3028;
   wire n_0_3029;
   wire n_0_3030;
   wire n_0_3031;
   wire n_0_3032;
   wire n_0_3033;
   wire n_0_3034;
   wire n_0_124_0;
   wire n_0_3036;
   wire n_0_3037;
   wire n_0_3035;
   wire n_0_125_0;
   wire n_0_125_1;
   wire n_0_125_2;
   wire n_0_125_3;
   wire n_0_125_4;
   wire n_0_125_5;
   wire n_0_125_6;
   wire n_0_125_7;
   wire n_0_125_8;
   wire n_0_125_9;
   wire n_0_125_10;
   wire n_0_125_11;
   wire n_0_125_12;
   wire n_0_125_13;
   wire n_0_125_14;
   wire n_0_125_15;
   wire n_0_125_16;
   wire n_0_125_17;
   wire n_0_125_18;
   wire n_0_125_19;
   wire n_0_125_20;
   wire n_0_125_21;
   wire n_0_125_22;
   wire n_0_125_23;
   wire n_0_125_24;
   wire n_0_125_25;
   wire n_0_125_26;
   wire n_0_125_27;
   wire n_0_125_28;
   wire n_0_125_29;
   wire n_0_125_30;
   wire n_0_125_31;
   wire n_0_125_32;

   assign product[63] = product[62];

   datapath i_0_0 (.multiplicand2(multiplicand2), .p_0({n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
      n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, uc_0}));
   AND2_X1 i_0_1_0 (.A1(multiplicand2[0]), .A2(multiplier2[0]), .ZN(product[0]));
   AND2_X1 i_0_1_1 (.A1(multiplier2[0]), .A2(n_0_0), .ZN(accumlator[1]));
   AND2_X1 i_0_1_2 (.A1(multiplier2[0]), .A2(n_0_1), .ZN(accumlator[2]));
   AND2_X1 i_0_1_3 (.A1(multiplier2[0]), .A2(n_0_2), .ZN(accumlator[3]));
   AND2_X1 i_0_1_4 (.A1(multiplier2[0]), .A2(n_0_3), .ZN(accumlator[4]));
   AND2_X1 i_0_1_5 (.A1(multiplier2[0]), .A2(n_0_4), .ZN(accumlator[5]));
   AND2_X1 i_0_1_6 (.A1(multiplier2[0]), .A2(n_0_5), .ZN(accumlator[6]));
   AND2_X1 i_0_1_7 (.A1(multiplier2[0]), .A2(n_0_6), .ZN(accumlator[7]));
   AND2_X1 i_0_1_8 (.A1(multiplier2[0]), .A2(n_0_7), .ZN(accumlator[8]));
   AND2_X1 i_0_1_9 (.A1(multiplier2[0]), .A2(n_0_8), .ZN(accumlator[9]));
   AND2_X1 i_0_1_10 (.A1(multiplier2[0]), .A2(n_0_9), .ZN(accumlator[10]));
   AND2_X1 i_0_1_11 (.A1(multiplier2[0]), .A2(n_0_10), .ZN(accumlator[11]));
   AND2_X1 i_0_1_12 (.A1(multiplier2[0]), .A2(n_0_11), .ZN(accumlator[12]));
   AND2_X1 i_0_1_13 (.A1(multiplier2[0]), .A2(n_0_12), .ZN(accumlator[13]));
   AND2_X1 i_0_1_14 (.A1(multiplier2[0]), .A2(n_0_13), .ZN(accumlator[14]));
   AND2_X1 i_0_1_15 (.A1(multiplier2[0]), .A2(n_0_14), .ZN(accumlator[15]));
   AND2_X1 i_0_1_16 (.A1(multiplier2[0]), .A2(n_0_15), .ZN(accumlator[16]));
   AND2_X1 i_0_1_17 (.A1(multiplier2[0]), .A2(n_0_16), .ZN(accumlator[17]));
   AND2_X1 i_0_1_18 (.A1(multiplier2[0]), .A2(n_0_17), .ZN(accumlator[18]));
   AND2_X1 i_0_1_19 (.A1(multiplier2[0]), .A2(n_0_18), .ZN(accumlator[19]));
   AND2_X1 i_0_1_20 (.A1(multiplier2[0]), .A2(n_0_19), .ZN(accumlator[20]));
   AND2_X1 i_0_1_21 (.A1(multiplier2[0]), .A2(n_0_20), .ZN(accumlator[21]));
   AND2_X1 i_0_1_22 (.A1(multiplier2[0]), .A2(n_0_21), .ZN(accumlator[22]));
   AND2_X1 i_0_1_23 (.A1(multiplier2[0]), .A2(n_0_22), .ZN(accumlator[23]));
   AND2_X1 i_0_1_24 (.A1(multiplier2[0]), .A2(n_0_23), .ZN(accumlator[24]));
   AND2_X1 i_0_1_25 (.A1(multiplier2[0]), .A2(n_0_24), .ZN(accumlator[25]));
   AND2_X1 i_0_1_26 (.A1(multiplier2[0]), .A2(n_0_25), .ZN(accumlator[26]));
   AND2_X1 i_0_1_27 (.A1(multiplier2[0]), .A2(n_0_26), .ZN(accumlator[27]));
   AND2_X1 i_0_1_28 (.A1(multiplier2[0]), .A2(n_0_27), .ZN(accumlator[28]));
   AND2_X1 i_0_1_29 (.A1(multiplier2[0]), .A2(n_0_28), .ZN(accumlator[29]));
   AND2_X1 i_0_1_30 (.A1(multiplier2[0]), .A2(n_0_29), .ZN(accumlator[30]));
   AND2_X1 i_0_1_31 (.A1(multiplier2[0]), .A2(n_0_30), .ZN(accumlator[31]));
   datapath__0_0 i_0_2 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_1, 
      accumlator[31], accumlator[30], accumlator[29], accumlator[28], 
      accumlator[27], accumlator[26], accumlator[25], accumlator[24], 
      accumlator[23], accumlator[22], accumlator[21], accumlator[20], 
      accumlator[19], accumlator[18], accumlator[17], accumlator[16], 
      accumlator[15], accumlator[14], accumlator[13], accumlator[12], 
      accumlator[11], accumlator[10], accumlator[9], accumlator[8], 
      accumlator[7], accumlator[6], accumlator[5], accumlator[4], accumlator[3], 
      accumlator[2], accumlator[1]}), .p_2({n_0_62, n_0_61, n_0_60, n_0_59, 
      n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, 
      n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, 
      n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, 
      n_0_31}));
   datapath__0_1 i_0_3 (.multiplicand2(multiplicand2), .p_0({uc_2, 
      accumlator[31], accumlator[30], accumlator[29], accumlator[28], 
      accumlator[27], accumlator[26], accumlator[25], accumlator[24], 
      accumlator[23], accumlator[22], accumlator[21], accumlator[20], 
      accumlator[19], accumlator[18], accumlator[17], accumlator[16], 
      accumlator[15], accumlator[14], accumlator[13], accumlator[12], 
      accumlator[11], accumlator[10], accumlator[9], accumlator[8], 
      accumlator[7], accumlator[6], accumlator[5], accumlator[4], accumlator[3], 
      accumlator[2], accumlator[1]}), .p_1({n_0_94, n_0_93, n_0_92, n_0_91, 
      n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, 
      n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, 
      n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, 
      n_0_63}));
   INV_X1 i_0_4_0 (.A(multiplier2[1]), .ZN(n_0_4_0));
   AND2_X1 i_0_4_1 (.A1(n_0_4_0), .A2(multiplier2[0]), .ZN(n_0_96));
   NOR2_X1 i_0_4_2 (.A1(n_0_4_0), .A2(multiplier2[0]), .ZN(n_0_97));
   NOR2_X1 i_0_4_3 (.A1(n_0_96), .A2(n_0_97), .ZN(n_0_95));
   AOI222_X1 i_0_5_0 (.A1(n_0_63), .A2(n_0_96), .B1(n_0_31), .B2(n_0_97), 
      .C1(accumlator[1]), .C2(n_0_95), .ZN(n_0_5_0));
   INV_X1 i_0_5_1 (.A(n_0_5_0), .ZN(product[1]));
   AOI222_X1 i_0_5_2 (.A1(n_0_96), .A2(n_0_64), .B1(n_0_97), .B2(n_0_32), 
      .C1(n_0_95), .C2(accumlator[2]), .ZN(n_0_5_1));
   INV_X1 i_0_5_3 (.A(n_0_5_1), .ZN(n_0_98));
   AOI222_X1 i_0_5_4 (.A1(n_0_96), .A2(n_0_65), .B1(n_0_97), .B2(n_0_33), 
      .C1(n_0_95), .C2(accumlator[3]), .ZN(n_0_5_2));
   INV_X1 i_0_5_5 (.A(n_0_5_2), .ZN(n_0_99));
   AOI222_X1 i_0_5_6 (.A1(n_0_96), .A2(n_0_66), .B1(n_0_97), .B2(n_0_34), 
      .C1(n_0_95), .C2(accumlator[4]), .ZN(n_0_5_3));
   INV_X1 i_0_5_7 (.A(n_0_5_3), .ZN(n_0_100));
   AOI222_X1 i_0_5_8 (.A1(n_0_96), .A2(n_0_67), .B1(n_0_97), .B2(n_0_35), 
      .C1(n_0_95), .C2(accumlator[5]), .ZN(n_0_5_4));
   INV_X1 i_0_5_9 (.A(n_0_5_4), .ZN(n_0_101));
   AOI222_X1 i_0_5_10 (.A1(n_0_96), .A2(n_0_68), .B1(n_0_97), .B2(n_0_36), 
      .C1(n_0_95), .C2(accumlator[6]), .ZN(n_0_5_5));
   INV_X1 i_0_5_11 (.A(n_0_5_5), .ZN(n_0_102));
   AOI222_X1 i_0_5_12 (.A1(n_0_96), .A2(n_0_69), .B1(n_0_97), .B2(n_0_37), 
      .C1(n_0_95), .C2(accumlator[7]), .ZN(n_0_5_6));
   INV_X1 i_0_5_13 (.A(n_0_5_6), .ZN(n_0_103));
   AOI222_X1 i_0_5_14 (.A1(n_0_96), .A2(n_0_70), .B1(n_0_97), .B2(n_0_38), 
      .C1(n_0_95), .C2(accumlator[8]), .ZN(n_0_5_7));
   INV_X1 i_0_5_15 (.A(n_0_5_7), .ZN(n_0_104));
   AOI222_X1 i_0_5_16 (.A1(n_0_96), .A2(n_0_71), .B1(n_0_97), .B2(n_0_39), 
      .C1(n_0_95), .C2(accumlator[9]), .ZN(n_0_5_8));
   INV_X1 i_0_5_17 (.A(n_0_5_8), .ZN(n_0_105));
   AOI222_X1 i_0_5_18 (.A1(n_0_96), .A2(n_0_72), .B1(n_0_97), .B2(n_0_40), 
      .C1(n_0_95), .C2(accumlator[10]), .ZN(n_0_5_9));
   INV_X1 i_0_5_19 (.A(n_0_5_9), .ZN(n_0_106));
   AOI222_X1 i_0_5_20 (.A1(n_0_96), .A2(n_0_73), .B1(n_0_97), .B2(n_0_41), 
      .C1(n_0_95), .C2(accumlator[11]), .ZN(n_0_5_10));
   INV_X1 i_0_5_21 (.A(n_0_5_10), .ZN(n_0_107));
   AOI222_X1 i_0_5_22 (.A1(n_0_96), .A2(n_0_74), .B1(n_0_97), .B2(n_0_42), 
      .C1(n_0_95), .C2(accumlator[12]), .ZN(n_0_5_11));
   INV_X1 i_0_5_23 (.A(n_0_5_11), .ZN(n_0_108));
   AOI222_X1 i_0_5_24 (.A1(n_0_96), .A2(n_0_75), .B1(n_0_97), .B2(n_0_43), 
      .C1(n_0_95), .C2(accumlator[13]), .ZN(n_0_5_12));
   INV_X1 i_0_5_25 (.A(n_0_5_12), .ZN(n_0_109));
   AOI222_X1 i_0_5_26 (.A1(n_0_96), .A2(n_0_76), .B1(n_0_97), .B2(n_0_44), 
      .C1(n_0_95), .C2(accumlator[14]), .ZN(n_0_5_13));
   INV_X1 i_0_5_27 (.A(n_0_5_13), .ZN(n_0_110));
   AOI222_X1 i_0_5_28 (.A1(n_0_96), .A2(n_0_77), .B1(n_0_97), .B2(n_0_45), 
      .C1(n_0_95), .C2(accumlator[15]), .ZN(n_0_5_14));
   INV_X1 i_0_5_29 (.A(n_0_5_14), .ZN(n_0_111));
   AOI222_X1 i_0_5_30 (.A1(n_0_96), .A2(n_0_78), .B1(n_0_97), .B2(n_0_46), 
      .C1(n_0_95), .C2(accumlator[16]), .ZN(n_0_5_15));
   INV_X1 i_0_5_31 (.A(n_0_5_15), .ZN(n_0_112));
   AOI222_X1 i_0_5_32 (.A1(n_0_96), .A2(n_0_79), .B1(n_0_97), .B2(n_0_47), 
      .C1(n_0_95), .C2(accumlator[17]), .ZN(n_0_5_16));
   INV_X1 i_0_5_33 (.A(n_0_5_16), .ZN(n_0_113));
   AOI222_X1 i_0_5_34 (.A1(n_0_96), .A2(n_0_80), .B1(n_0_97), .B2(n_0_48), 
      .C1(n_0_95), .C2(accumlator[18]), .ZN(n_0_5_17));
   INV_X1 i_0_5_35 (.A(n_0_5_17), .ZN(n_0_114));
   AOI222_X1 i_0_5_36 (.A1(n_0_96), .A2(n_0_81), .B1(n_0_97), .B2(n_0_49), 
      .C1(n_0_95), .C2(accumlator[19]), .ZN(n_0_5_18));
   INV_X1 i_0_5_37 (.A(n_0_5_18), .ZN(n_0_115));
   AOI222_X1 i_0_5_38 (.A1(n_0_96), .A2(n_0_82), .B1(n_0_97), .B2(n_0_50), 
      .C1(n_0_95), .C2(accumlator[20]), .ZN(n_0_5_19));
   INV_X1 i_0_5_39 (.A(n_0_5_19), .ZN(n_0_116));
   AOI222_X1 i_0_5_40 (.A1(n_0_96), .A2(n_0_83), .B1(n_0_97), .B2(n_0_51), 
      .C1(n_0_95), .C2(accumlator[21]), .ZN(n_0_5_20));
   INV_X1 i_0_5_41 (.A(n_0_5_20), .ZN(n_0_117));
   AOI222_X1 i_0_5_42 (.A1(n_0_96), .A2(n_0_84), .B1(n_0_97), .B2(n_0_52), 
      .C1(n_0_95), .C2(accumlator[22]), .ZN(n_0_5_21));
   INV_X1 i_0_5_43 (.A(n_0_5_21), .ZN(n_0_118));
   AOI222_X1 i_0_5_44 (.A1(n_0_96), .A2(n_0_85), .B1(n_0_97), .B2(n_0_53), 
      .C1(n_0_95), .C2(accumlator[23]), .ZN(n_0_5_22));
   INV_X1 i_0_5_45 (.A(n_0_5_22), .ZN(n_0_119));
   AOI222_X1 i_0_5_46 (.A1(n_0_96), .A2(n_0_86), .B1(n_0_97), .B2(n_0_54), 
      .C1(n_0_95), .C2(accumlator[24]), .ZN(n_0_5_23));
   INV_X1 i_0_5_47 (.A(n_0_5_23), .ZN(n_0_120));
   AOI222_X1 i_0_5_48 (.A1(n_0_96), .A2(n_0_87), .B1(n_0_97), .B2(n_0_55), 
      .C1(n_0_95), .C2(accumlator[25]), .ZN(n_0_5_24));
   INV_X1 i_0_5_49 (.A(n_0_5_24), .ZN(n_0_121));
   AOI222_X1 i_0_5_50 (.A1(n_0_96), .A2(n_0_88), .B1(n_0_97), .B2(n_0_56), 
      .C1(n_0_95), .C2(accumlator[26]), .ZN(n_0_5_25));
   INV_X1 i_0_5_51 (.A(n_0_5_25), .ZN(n_0_122));
   AOI222_X1 i_0_5_52 (.A1(n_0_96), .A2(n_0_89), .B1(n_0_97), .B2(n_0_57), 
      .C1(n_0_95), .C2(accumlator[27]), .ZN(n_0_5_26));
   INV_X1 i_0_5_53 (.A(n_0_5_26), .ZN(n_0_123));
   AOI222_X1 i_0_5_54 (.A1(n_0_96), .A2(n_0_90), .B1(n_0_97), .B2(n_0_58), 
      .C1(n_0_95), .C2(accumlator[28]), .ZN(n_0_5_27));
   INV_X1 i_0_5_55 (.A(n_0_5_27), .ZN(n_0_124));
   AOI222_X1 i_0_5_56 (.A1(n_0_96), .A2(n_0_91), .B1(n_0_97), .B2(n_0_59), 
      .C1(n_0_95), .C2(accumlator[29]), .ZN(n_0_5_28));
   INV_X1 i_0_5_57 (.A(n_0_5_28), .ZN(n_0_125));
   AOI222_X1 i_0_5_58 (.A1(n_0_96), .A2(n_0_92), .B1(n_0_97), .B2(n_0_60), 
      .C1(n_0_95), .C2(accumlator[30]), .ZN(n_0_5_29));
   INV_X1 i_0_5_59 (.A(n_0_5_29), .ZN(n_0_126));
   AND2_X1 i_0_5_60 (.A1(n_0_95), .A2(accumlator[31]), .ZN(n_0_5_30));
   AOI221_X1 i_0_5_61 (.A(n_0_5_30), .B1(n_0_96), .B2(n_0_93), .C1(n_0_97), 
      .C2(n_0_61), .ZN(n_0_5_31));
   INV_X1 i_0_5_62 (.A(n_0_5_31), .ZN(n_0_127));
   AOI221_X1 i_0_5_63 (.A(n_0_5_30), .B1(n_0_96), .B2(n_0_94), .C1(n_0_97), 
      .C2(n_0_62), .ZN(n_0_5_32));
   INV_X1 i_0_5_64 (.A(n_0_5_32), .ZN(n_0_128));
   datapath__0_4 i_0_6 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_3, 
      n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
      n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, 
      n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, 
      n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98}), .p_2({
      n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, 
      n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, 
      n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, 
      n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129}));
   datapath__0_5 i_0_7 (.multiplicand2(multiplicand2), .p_0({uc_4, n_0_128, 
      n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98}), .p_1({n_0_192, 
      n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, 
      n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, 
      n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, 
      n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161}));
   INV_X1 i_0_8_0 (.A(multiplier2[2]), .ZN(n_0_8_0));
   AND2_X1 i_0_8_1 (.A1(n_0_8_0), .A2(multiplier2[1]), .ZN(n_0_194));
   NOR2_X1 i_0_8_2 (.A1(n_0_8_0), .A2(multiplier2[1]), .ZN(n_0_195));
   NOR2_X1 i_0_8_3 (.A1(n_0_194), .A2(n_0_195), .ZN(n_0_193));
   AOI222_X1 i_0_9_0 (.A1(n_0_161), .A2(n_0_194), .B1(n_0_129), .B2(n_0_195), 
      .C1(n_0_98), .C2(n_0_193), .ZN(n_0_9_0));
   INV_X1 i_0_9_1 (.A(n_0_9_0), .ZN(product[2]));
   AOI222_X1 i_0_9_2 (.A1(n_0_194), .A2(n_0_162), .B1(n_0_195), .B2(n_0_130), 
      .C1(n_0_193), .C2(n_0_99), .ZN(n_0_9_1));
   INV_X1 i_0_9_3 (.A(n_0_9_1), .ZN(n_0_196));
   AOI222_X1 i_0_9_4 (.A1(n_0_194), .A2(n_0_163), .B1(n_0_195), .B2(n_0_131), 
      .C1(n_0_193), .C2(n_0_100), .ZN(n_0_9_2));
   INV_X1 i_0_9_5 (.A(n_0_9_2), .ZN(n_0_197));
   AOI222_X1 i_0_9_6 (.A1(n_0_194), .A2(n_0_164), .B1(n_0_195), .B2(n_0_132), 
      .C1(n_0_193), .C2(n_0_101), .ZN(n_0_9_3));
   INV_X1 i_0_9_7 (.A(n_0_9_3), .ZN(n_0_198));
   AOI222_X1 i_0_9_8 (.A1(n_0_194), .A2(n_0_165), .B1(n_0_195), .B2(n_0_133), 
      .C1(n_0_193), .C2(n_0_102), .ZN(n_0_9_4));
   INV_X1 i_0_9_9 (.A(n_0_9_4), .ZN(n_0_199));
   AOI222_X1 i_0_9_10 (.A1(n_0_194), .A2(n_0_166), .B1(n_0_195), .B2(n_0_134), 
      .C1(n_0_193), .C2(n_0_103), .ZN(n_0_9_5));
   INV_X1 i_0_9_11 (.A(n_0_9_5), .ZN(n_0_200));
   AOI222_X1 i_0_9_12 (.A1(n_0_194), .A2(n_0_167), .B1(n_0_195), .B2(n_0_135), 
      .C1(n_0_193), .C2(n_0_104), .ZN(n_0_9_6));
   INV_X1 i_0_9_13 (.A(n_0_9_6), .ZN(n_0_201));
   AOI222_X1 i_0_9_14 (.A1(n_0_194), .A2(n_0_168), .B1(n_0_195), .B2(n_0_136), 
      .C1(n_0_193), .C2(n_0_105), .ZN(n_0_9_7));
   INV_X1 i_0_9_15 (.A(n_0_9_7), .ZN(n_0_202));
   AOI222_X1 i_0_9_16 (.A1(n_0_194), .A2(n_0_169), .B1(n_0_195), .B2(n_0_137), 
      .C1(n_0_193), .C2(n_0_106), .ZN(n_0_9_8));
   INV_X1 i_0_9_17 (.A(n_0_9_8), .ZN(n_0_203));
   AOI222_X1 i_0_9_18 (.A1(n_0_194), .A2(n_0_170), .B1(n_0_195), .B2(n_0_138), 
      .C1(n_0_193), .C2(n_0_107), .ZN(n_0_9_9));
   INV_X1 i_0_9_19 (.A(n_0_9_9), .ZN(n_0_204));
   AOI222_X1 i_0_9_20 (.A1(n_0_194), .A2(n_0_171), .B1(n_0_195), .B2(n_0_139), 
      .C1(n_0_193), .C2(n_0_108), .ZN(n_0_9_10));
   INV_X1 i_0_9_21 (.A(n_0_9_10), .ZN(n_0_205));
   AOI222_X1 i_0_9_22 (.A1(n_0_194), .A2(n_0_172), .B1(n_0_195), .B2(n_0_140), 
      .C1(n_0_193), .C2(n_0_109), .ZN(n_0_9_11));
   INV_X1 i_0_9_23 (.A(n_0_9_11), .ZN(n_0_206));
   AOI222_X1 i_0_9_24 (.A1(n_0_194), .A2(n_0_173), .B1(n_0_195), .B2(n_0_141), 
      .C1(n_0_193), .C2(n_0_110), .ZN(n_0_9_12));
   INV_X1 i_0_9_25 (.A(n_0_9_12), .ZN(n_0_207));
   AOI222_X1 i_0_9_26 (.A1(n_0_194), .A2(n_0_174), .B1(n_0_195), .B2(n_0_142), 
      .C1(n_0_193), .C2(n_0_111), .ZN(n_0_9_13));
   INV_X1 i_0_9_27 (.A(n_0_9_13), .ZN(n_0_208));
   AOI222_X1 i_0_9_28 (.A1(n_0_194), .A2(n_0_175), .B1(n_0_195), .B2(n_0_143), 
      .C1(n_0_193), .C2(n_0_112), .ZN(n_0_9_14));
   INV_X1 i_0_9_29 (.A(n_0_9_14), .ZN(n_0_209));
   AOI222_X1 i_0_9_30 (.A1(n_0_194), .A2(n_0_176), .B1(n_0_195), .B2(n_0_144), 
      .C1(n_0_193), .C2(n_0_113), .ZN(n_0_9_15));
   INV_X1 i_0_9_31 (.A(n_0_9_15), .ZN(n_0_210));
   AOI222_X1 i_0_9_32 (.A1(n_0_194), .A2(n_0_177), .B1(n_0_195), .B2(n_0_145), 
      .C1(n_0_193), .C2(n_0_114), .ZN(n_0_9_16));
   INV_X1 i_0_9_33 (.A(n_0_9_16), .ZN(n_0_211));
   AOI222_X1 i_0_9_34 (.A1(n_0_194), .A2(n_0_178), .B1(n_0_195), .B2(n_0_146), 
      .C1(n_0_193), .C2(n_0_115), .ZN(n_0_9_17));
   INV_X1 i_0_9_35 (.A(n_0_9_17), .ZN(n_0_212));
   AOI222_X1 i_0_9_36 (.A1(n_0_194), .A2(n_0_179), .B1(n_0_195), .B2(n_0_147), 
      .C1(n_0_193), .C2(n_0_116), .ZN(n_0_9_18));
   INV_X1 i_0_9_37 (.A(n_0_9_18), .ZN(n_0_213));
   AOI222_X1 i_0_9_38 (.A1(n_0_194), .A2(n_0_180), .B1(n_0_195), .B2(n_0_148), 
      .C1(n_0_193), .C2(n_0_117), .ZN(n_0_9_19));
   INV_X1 i_0_9_39 (.A(n_0_9_19), .ZN(n_0_214));
   AOI222_X1 i_0_9_40 (.A1(n_0_194), .A2(n_0_181), .B1(n_0_195), .B2(n_0_149), 
      .C1(n_0_193), .C2(n_0_118), .ZN(n_0_9_20));
   INV_X1 i_0_9_41 (.A(n_0_9_20), .ZN(n_0_215));
   AOI222_X1 i_0_9_42 (.A1(n_0_194), .A2(n_0_182), .B1(n_0_195), .B2(n_0_150), 
      .C1(n_0_193), .C2(n_0_119), .ZN(n_0_9_21));
   INV_X1 i_0_9_43 (.A(n_0_9_21), .ZN(n_0_216));
   AOI222_X1 i_0_9_44 (.A1(n_0_194), .A2(n_0_183), .B1(n_0_195), .B2(n_0_151), 
      .C1(n_0_193), .C2(n_0_120), .ZN(n_0_9_22));
   INV_X1 i_0_9_45 (.A(n_0_9_22), .ZN(n_0_217));
   AOI222_X1 i_0_9_46 (.A1(n_0_194), .A2(n_0_184), .B1(n_0_195), .B2(n_0_152), 
      .C1(n_0_193), .C2(n_0_121), .ZN(n_0_9_23));
   INV_X1 i_0_9_47 (.A(n_0_9_23), .ZN(n_0_218));
   AOI222_X1 i_0_9_48 (.A1(n_0_194), .A2(n_0_185), .B1(n_0_195), .B2(n_0_153), 
      .C1(n_0_193), .C2(n_0_122), .ZN(n_0_9_24));
   INV_X1 i_0_9_49 (.A(n_0_9_24), .ZN(n_0_219));
   AOI222_X1 i_0_9_50 (.A1(n_0_194), .A2(n_0_186), .B1(n_0_195), .B2(n_0_154), 
      .C1(n_0_193), .C2(n_0_123), .ZN(n_0_9_25));
   INV_X1 i_0_9_51 (.A(n_0_9_25), .ZN(n_0_220));
   AOI222_X1 i_0_9_52 (.A1(n_0_194), .A2(n_0_187), .B1(n_0_195), .B2(n_0_155), 
      .C1(n_0_193), .C2(n_0_124), .ZN(n_0_9_26));
   INV_X1 i_0_9_53 (.A(n_0_9_26), .ZN(n_0_221));
   AOI222_X1 i_0_9_54 (.A1(n_0_194), .A2(n_0_188), .B1(n_0_195), .B2(n_0_156), 
      .C1(n_0_193), .C2(n_0_125), .ZN(n_0_9_27));
   INV_X1 i_0_9_55 (.A(n_0_9_27), .ZN(n_0_222));
   AOI222_X1 i_0_9_56 (.A1(n_0_194), .A2(n_0_189), .B1(n_0_195), .B2(n_0_157), 
      .C1(n_0_193), .C2(n_0_126), .ZN(n_0_9_28));
   INV_X1 i_0_9_57 (.A(n_0_9_28), .ZN(n_0_223));
   AOI222_X1 i_0_9_58 (.A1(n_0_194), .A2(n_0_190), .B1(n_0_195), .B2(n_0_158), 
      .C1(n_0_193), .C2(n_0_127), .ZN(n_0_9_29));
   INV_X1 i_0_9_59 (.A(n_0_9_29), .ZN(n_0_224));
   AND2_X1 i_0_9_60 (.A1(n_0_193), .A2(n_0_128), .ZN(n_0_9_30));
   AOI221_X1 i_0_9_61 (.A(n_0_9_30), .B1(n_0_194), .B2(n_0_191), .C1(n_0_195), 
      .C2(n_0_159), .ZN(n_0_9_31));
   INV_X1 i_0_9_62 (.A(n_0_9_31), .ZN(n_0_225));
   AOI221_X1 i_0_9_63 (.A(n_0_9_30), .B1(n_0_194), .B2(n_0_192), .C1(n_0_195), 
      .C2(n_0_160), .ZN(n_0_9_32));
   INV_X1 i_0_9_64 (.A(n_0_9_32), .ZN(n_0_226));
   datapath__0_8 i_0_10 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_5, 
      n_0_226, n_0_225, n_0_224, n_0_223, n_0_222, n_0_221, n_0_220, n_0_219, 
      n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, 
      n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, 
      n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196}), .p_2({
      n_0_258, n_0_257, n_0_256, n_0_255, n_0_254, n_0_253, n_0_252, n_0_251, 
      n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, 
      n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, 
      n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, n_0_229, n_0_228, n_0_227}));
   datapath__0_9 i_0_11 (.multiplicand2(multiplicand2), .p_0({uc_6, n_0_226, 
      n_0_225, n_0_224, n_0_223, n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, 
      n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, 
      n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, 
      n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196}), .p_1({n_0_290, 
      n_0_289, n_0_288, n_0_287, n_0_286, n_0_285, n_0_284, n_0_283, n_0_282, 
      n_0_281, n_0_280, n_0_279, n_0_278, n_0_277, n_0_276, n_0_275, n_0_274, 
      n_0_273, n_0_272, n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, n_0_266, 
      n_0_265, n_0_264, n_0_263, n_0_262, n_0_261, n_0_260, n_0_259}));
   INV_X1 i_0_12_0 (.A(multiplier2[3]), .ZN(n_0_12_0));
   AND2_X1 i_0_12_1 (.A1(n_0_12_0), .A2(multiplier2[2]), .ZN(n_0_292));
   NOR2_X1 i_0_12_2 (.A1(n_0_12_0), .A2(multiplier2[2]), .ZN(n_0_293));
   NOR2_X1 i_0_12_3 (.A1(n_0_292), .A2(n_0_293), .ZN(n_0_291));
   AOI222_X1 i_0_13_0 (.A1(n_0_259), .A2(n_0_292), .B1(n_0_227), .B2(n_0_293), 
      .C1(n_0_196), .C2(n_0_291), .ZN(n_0_13_0));
   INV_X1 i_0_13_1 (.A(n_0_13_0), .ZN(product[3]));
   AOI222_X1 i_0_13_2 (.A1(n_0_292), .A2(n_0_260), .B1(n_0_293), .B2(n_0_228), 
      .C1(n_0_291), .C2(n_0_197), .ZN(n_0_13_1));
   INV_X1 i_0_13_3 (.A(n_0_13_1), .ZN(n_0_294));
   AOI222_X1 i_0_13_4 (.A1(n_0_292), .A2(n_0_261), .B1(n_0_293), .B2(n_0_229), 
      .C1(n_0_291), .C2(n_0_198), .ZN(n_0_13_2));
   INV_X1 i_0_13_5 (.A(n_0_13_2), .ZN(n_0_295));
   AOI222_X1 i_0_13_6 (.A1(n_0_292), .A2(n_0_262), .B1(n_0_293), .B2(n_0_230), 
      .C1(n_0_291), .C2(n_0_199), .ZN(n_0_13_3));
   INV_X1 i_0_13_7 (.A(n_0_13_3), .ZN(n_0_296));
   AOI222_X1 i_0_13_8 (.A1(n_0_292), .A2(n_0_263), .B1(n_0_293), .B2(n_0_231), 
      .C1(n_0_291), .C2(n_0_200), .ZN(n_0_13_4));
   INV_X1 i_0_13_9 (.A(n_0_13_4), .ZN(n_0_297));
   AOI222_X1 i_0_13_10 (.A1(n_0_292), .A2(n_0_264), .B1(n_0_293), .B2(n_0_232), 
      .C1(n_0_291), .C2(n_0_201), .ZN(n_0_13_5));
   INV_X1 i_0_13_11 (.A(n_0_13_5), .ZN(n_0_298));
   AOI222_X1 i_0_13_12 (.A1(n_0_292), .A2(n_0_265), .B1(n_0_293), .B2(n_0_233), 
      .C1(n_0_291), .C2(n_0_202), .ZN(n_0_13_6));
   INV_X1 i_0_13_13 (.A(n_0_13_6), .ZN(n_0_299));
   AOI222_X1 i_0_13_14 (.A1(n_0_292), .A2(n_0_266), .B1(n_0_293), .B2(n_0_234), 
      .C1(n_0_291), .C2(n_0_203), .ZN(n_0_13_7));
   INV_X1 i_0_13_15 (.A(n_0_13_7), .ZN(n_0_300));
   AOI222_X1 i_0_13_16 (.A1(n_0_292), .A2(n_0_267), .B1(n_0_293), .B2(n_0_235), 
      .C1(n_0_291), .C2(n_0_204), .ZN(n_0_13_8));
   INV_X1 i_0_13_17 (.A(n_0_13_8), .ZN(n_0_301));
   AOI222_X1 i_0_13_18 (.A1(n_0_292), .A2(n_0_268), .B1(n_0_293), .B2(n_0_236), 
      .C1(n_0_291), .C2(n_0_205), .ZN(n_0_13_9));
   INV_X1 i_0_13_19 (.A(n_0_13_9), .ZN(n_0_302));
   AOI222_X1 i_0_13_20 (.A1(n_0_292), .A2(n_0_269), .B1(n_0_293), .B2(n_0_237), 
      .C1(n_0_291), .C2(n_0_206), .ZN(n_0_13_10));
   INV_X1 i_0_13_21 (.A(n_0_13_10), .ZN(n_0_303));
   AOI222_X1 i_0_13_22 (.A1(n_0_292), .A2(n_0_270), .B1(n_0_293), .B2(n_0_238), 
      .C1(n_0_291), .C2(n_0_207), .ZN(n_0_13_11));
   INV_X1 i_0_13_23 (.A(n_0_13_11), .ZN(n_0_304));
   AOI222_X1 i_0_13_24 (.A1(n_0_292), .A2(n_0_271), .B1(n_0_293), .B2(n_0_239), 
      .C1(n_0_291), .C2(n_0_208), .ZN(n_0_13_12));
   INV_X1 i_0_13_25 (.A(n_0_13_12), .ZN(n_0_305));
   AOI222_X1 i_0_13_26 (.A1(n_0_292), .A2(n_0_272), .B1(n_0_293), .B2(n_0_240), 
      .C1(n_0_291), .C2(n_0_209), .ZN(n_0_13_13));
   INV_X1 i_0_13_27 (.A(n_0_13_13), .ZN(n_0_306));
   AOI222_X1 i_0_13_28 (.A1(n_0_292), .A2(n_0_273), .B1(n_0_293), .B2(n_0_241), 
      .C1(n_0_291), .C2(n_0_210), .ZN(n_0_13_14));
   INV_X1 i_0_13_29 (.A(n_0_13_14), .ZN(n_0_307));
   AOI222_X1 i_0_13_30 (.A1(n_0_292), .A2(n_0_274), .B1(n_0_293), .B2(n_0_242), 
      .C1(n_0_291), .C2(n_0_211), .ZN(n_0_13_15));
   INV_X1 i_0_13_31 (.A(n_0_13_15), .ZN(n_0_308));
   AOI222_X1 i_0_13_32 (.A1(n_0_292), .A2(n_0_275), .B1(n_0_293), .B2(n_0_243), 
      .C1(n_0_291), .C2(n_0_212), .ZN(n_0_13_16));
   INV_X1 i_0_13_33 (.A(n_0_13_16), .ZN(n_0_309));
   AOI222_X1 i_0_13_34 (.A1(n_0_292), .A2(n_0_276), .B1(n_0_293), .B2(n_0_244), 
      .C1(n_0_291), .C2(n_0_213), .ZN(n_0_13_17));
   INV_X1 i_0_13_35 (.A(n_0_13_17), .ZN(n_0_310));
   AOI222_X1 i_0_13_36 (.A1(n_0_292), .A2(n_0_277), .B1(n_0_293), .B2(n_0_245), 
      .C1(n_0_291), .C2(n_0_214), .ZN(n_0_13_18));
   INV_X1 i_0_13_37 (.A(n_0_13_18), .ZN(n_0_311));
   AOI222_X1 i_0_13_38 (.A1(n_0_292), .A2(n_0_278), .B1(n_0_293), .B2(n_0_246), 
      .C1(n_0_291), .C2(n_0_215), .ZN(n_0_13_19));
   INV_X1 i_0_13_39 (.A(n_0_13_19), .ZN(n_0_312));
   AOI222_X1 i_0_13_40 (.A1(n_0_292), .A2(n_0_279), .B1(n_0_293), .B2(n_0_247), 
      .C1(n_0_291), .C2(n_0_216), .ZN(n_0_13_20));
   INV_X1 i_0_13_41 (.A(n_0_13_20), .ZN(n_0_313));
   AOI222_X1 i_0_13_42 (.A1(n_0_292), .A2(n_0_280), .B1(n_0_293), .B2(n_0_248), 
      .C1(n_0_291), .C2(n_0_217), .ZN(n_0_13_21));
   INV_X1 i_0_13_43 (.A(n_0_13_21), .ZN(n_0_314));
   AOI222_X1 i_0_13_44 (.A1(n_0_292), .A2(n_0_281), .B1(n_0_293), .B2(n_0_249), 
      .C1(n_0_291), .C2(n_0_218), .ZN(n_0_13_22));
   INV_X1 i_0_13_45 (.A(n_0_13_22), .ZN(n_0_315));
   AOI222_X1 i_0_13_46 (.A1(n_0_292), .A2(n_0_282), .B1(n_0_293), .B2(n_0_250), 
      .C1(n_0_291), .C2(n_0_219), .ZN(n_0_13_23));
   INV_X1 i_0_13_47 (.A(n_0_13_23), .ZN(n_0_316));
   AOI222_X1 i_0_13_48 (.A1(n_0_292), .A2(n_0_283), .B1(n_0_293), .B2(n_0_251), 
      .C1(n_0_291), .C2(n_0_220), .ZN(n_0_13_24));
   INV_X1 i_0_13_49 (.A(n_0_13_24), .ZN(n_0_317));
   AOI222_X1 i_0_13_50 (.A1(n_0_292), .A2(n_0_284), .B1(n_0_293), .B2(n_0_252), 
      .C1(n_0_291), .C2(n_0_221), .ZN(n_0_13_25));
   INV_X1 i_0_13_51 (.A(n_0_13_25), .ZN(n_0_318));
   AOI222_X1 i_0_13_52 (.A1(n_0_292), .A2(n_0_285), .B1(n_0_293), .B2(n_0_253), 
      .C1(n_0_291), .C2(n_0_222), .ZN(n_0_13_26));
   INV_X1 i_0_13_53 (.A(n_0_13_26), .ZN(n_0_319));
   AOI222_X1 i_0_13_54 (.A1(n_0_292), .A2(n_0_286), .B1(n_0_293), .B2(n_0_254), 
      .C1(n_0_291), .C2(n_0_223), .ZN(n_0_13_27));
   INV_X1 i_0_13_55 (.A(n_0_13_27), .ZN(n_0_320));
   AOI222_X1 i_0_13_56 (.A1(n_0_292), .A2(n_0_287), .B1(n_0_293), .B2(n_0_255), 
      .C1(n_0_291), .C2(n_0_224), .ZN(n_0_13_28));
   INV_X1 i_0_13_57 (.A(n_0_13_28), .ZN(n_0_321));
   AOI222_X1 i_0_13_58 (.A1(n_0_292), .A2(n_0_288), .B1(n_0_293), .B2(n_0_256), 
      .C1(n_0_291), .C2(n_0_225), .ZN(n_0_13_29));
   INV_X1 i_0_13_59 (.A(n_0_13_29), .ZN(n_0_322));
   AND2_X1 i_0_13_60 (.A1(n_0_291), .A2(n_0_226), .ZN(n_0_13_30));
   AOI221_X1 i_0_13_61 (.A(n_0_13_30), .B1(n_0_292), .B2(n_0_289), .C1(n_0_293), 
      .C2(n_0_257), .ZN(n_0_13_31));
   INV_X1 i_0_13_62 (.A(n_0_13_31), .ZN(n_0_323));
   AOI221_X1 i_0_13_63 (.A(n_0_13_30), .B1(n_0_292), .B2(n_0_290), .C1(n_0_293), 
      .C2(n_0_258), .ZN(n_0_13_32));
   INV_X1 i_0_13_64 (.A(n_0_13_32), .ZN(n_0_324));
   datapath__0_12 i_0_14 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_7, 
      n_0_324, n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, 
      n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, n_0_309, 
      n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, n_0_302, n_0_301, 
      n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, n_0_294}), .p_2({
      n_0_356, n_0_355, n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, n_0_349, 
      n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, n_0_342, n_0_341, 
      n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, 
      n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325}));
   datapath__0_13 i_0_15 (.multiplicand2(multiplicand2), .p_0({uc_8, n_0_324, 
      n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, 
      n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, n_0_309, n_0_308, 
      n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, n_0_302, n_0_301, n_0_300, 
      n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, n_0_294}), .p_1({n_0_388, 
      n_0_387, n_0_386, n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, 
      n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, 
      n_0_371, n_0_370, n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, n_0_364, 
      n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357}));
   INV_X1 i_0_16_0 (.A(multiplier2[4]), .ZN(n_0_16_0));
   AND2_X1 i_0_16_1 (.A1(n_0_16_0), .A2(multiplier2[3]), .ZN(n_0_390));
   NOR2_X1 i_0_16_2 (.A1(n_0_16_0), .A2(multiplier2[3]), .ZN(n_0_391));
   NOR2_X1 i_0_16_3 (.A1(n_0_390), .A2(n_0_391), .ZN(n_0_389));
   AOI222_X1 i_0_17_0 (.A1(n_0_357), .A2(n_0_390), .B1(n_0_325), .B2(n_0_391), 
      .C1(n_0_294), .C2(n_0_389), .ZN(n_0_17_0));
   INV_X1 i_0_17_1 (.A(n_0_17_0), .ZN(product[4]));
   AOI222_X1 i_0_17_2 (.A1(n_0_390), .A2(n_0_358), .B1(n_0_391), .B2(n_0_326), 
      .C1(n_0_389), .C2(n_0_295), .ZN(n_0_17_1));
   INV_X1 i_0_17_3 (.A(n_0_17_1), .ZN(n_0_392));
   AOI222_X1 i_0_17_4 (.A1(n_0_390), .A2(n_0_359), .B1(n_0_391), .B2(n_0_327), 
      .C1(n_0_389), .C2(n_0_296), .ZN(n_0_17_2));
   INV_X1 i_0_17_5 (.A(n_0_17_2), .ZN(n_0_393));
   AOI222_X1 i_0_17_6 (.A1(n_0_390), .A2(n_0_360), .B1(n_0_391), .B2(n_0_328), 
      .C1(n_0_389), .C2(n_0_297), .ZN(n_0_17_3));
   INV_X1 i_0_17_7 (.A(n_0_17_3), .ZN(n_0_394));
   AOI222_X1 i_0_17_8 (.A1(n_0_390), .A2(n_0_361), .B1(n_0_391), .B2(n_0_329), 
      .C1(n_0_389), .C2(n_0_298), .ZN(n_0_17_4));
   INV_X1 i_0_17_9 (.A(n_0_17_4), .ZN(n_0_395));
   AOI222_X1 i_0_17_10 (.A1(n_0_390), .A2(n_0_362), .B1(n_0_391), .B2(n_0_330), 
      .C1(n_0_389), .C2(n_0_299), .ZN(n_0_17_5));
   INV_X1 i_0_17_11 (.A(n_0_17_5), .ZN(n_0_396));
   AOI222_X1 i_0_17_12 (.A1(n_0_390), .A2(n_0_363), .B1(n_0_391), .B2(n_0_331), 
      .C1(n_0_389), .C2(n_0_300), .ZN(n_0_17_6));
   INV_X1 i_0_17_13 (.A(n_0_17_6), .ZN(n_0_397));
   AOI222_X1 i_0_17_14 (.A1(n_0_390), .A2(n_0_364), .B1(n_0_391), .B2(n_0_332), 
      .C1(n_0_389), .C2(n_0_301), .ZN(n_0_17_7));
   INV_X1 i_0_17_15 (.A(n_0_17_7), .ZN(n_0_398));
   AOI222_X1 i_0_17_16 (.A1(n_0_390), .A2(n_0_365), .B1(n_0_391), .B2(n_0_333), 
      .C1(n_0_389), .C2(n_0_302), .ZN(n_0_17_8));
   INV_X1 i_0_17_17 (.A(n_0_17_8), .ZN(n_0_399));
   AOI222_X1 i_0_17_18 (.A1(n_0_390), .A2(n_0_366), .B1(n_0_391), .B2(n_0_334), 
      .C1(n_0_389), .C2(n_0_303), .ZN(n_0_17_9));
   INV_X1 i_0_17_19 (.A(n_0_17_9), .ZN(n_0_400));
   AOI222_X1 i_0_17_20 (.A1(n_0_390), .A2(n_0_367), .B1(n_0_391), .B2(n_0_335), 
      .C1(n_0_389), .C2(n_0_304), .ZN(n_0_17_10));
   INV_X1 i_0_17_21 (.A(n_0_17_10), .ZN(n_0_401));
   AOI222_X1 i_0_17_22 (.A1(n_0_390), .A2(n_0_368), .B1(n_0_391), .B2(n_0_336), 
      .C1(n_0_389), .C2(n_0_305), .ZN(n_0_17_11));
   INV_X1 i_0_17_23 (.A(n_0_17_11), .ZN(n_0_402));
   AOI222_X1 i_0_17_24 (.A1(n_0_390), .A2(n_0_369), .B1(n_0_391), .B2(n_0_337), 
      .C1(n_0_389), .C2(n_0_306), .ZN(n_0_17_12));
   INV_X1 i_0_17_25 (.A(n_0_17_12), .ZN(n_0_403));
   AOI222_X1 i_0_17_26 (.A1(n_0_390), .A2(n_0_370), .B1(n_0_391), .B2(n_0_338), 
      .C1(n_0_389), .C2(n_0_307), .ZN(n_0_17_13));
   INV_X1 i_0_17_27 (.A(n_0_17_13), .ZN(n_0_404));
   AOI222_X1 i_0_17_28 (.A1(n_0_390), .A2(n_0_371), .B1(n_0_391), .B2(n_0_339), 
      .C1(n_0_389), .C2(n_0_308), .ZN(n_0_17_14));
   INV_X1 i_0_17_29 (.A(n_0_17_14), .ZN(n_0_405));
   AOI222_X1 i_0_17_30 (.A1(n_0_390), .A2(n_0_372), .B1(n_0_391), .B2(n_0_340), 
      .C1(n_0_389), .C2(n_0_309), .ZN(n_0_17_15));
   INV_X1 i_0_17_31 (.A(n_0_17_15), .ZN(n_0_406));
   AOI222_X1 i_0_17_32 (.A1(n_0_390), .A2(n_0_373), .B1(n_0_391), .B2(n_0_341), 
      .C1(n_0_389), .C2(n_0_310), .ZN(n_0_17_16));
   INV_X1 i_0_17_33 (.A(n_0_17_16), .ZN(n_0_407));
   AOI222_X1 i_0_17_34 (.A1(n_0_390), .A2(n_0_374), .B1(n_0_391), .B2(n_0_342), 
      .C1(n_0_389), .C2(n_0_311), .ZN(n_0_17_17));
   INV_X1 i_0_17_35 (.A(n_0_17_17), .ZN(n_0_408));
   AOI222_X1 i_0_17_36 (.A1(n_0_390), .A2(n_0_375), .B1(n_0_391), .B2(n_0_343), 
      .C1(n_0_389), .C2(n_0_312), .ZN(n_0_17_18));
   INV_X1 i_0_17_37 (.A(n_0_17_18), .ZN(n_0_409));
   AOI222_X1 i_0_17_38 (.A1(n_0_390), .A2(n_0_376), .B1(n_0_391), .B2(n_0_344), 
      .C1(n_0_389), .C2(n_0_313), .ZN(n_0_17_19));
   INV_X1 i_0_17_39 (.A(n_0_17_19), .ZN(n_0_410));
   AOI222_X1 i_0_17_40 (.A1(n_0_390), .A2(n_0_377), .B1(n_0_391), .B2(n_0_345), 
      .C1(n_0_389), .C2(n_0_314), .ZN(n_0_17_20));
   INV_X1 i_0_17_41 (.A(n_0_17_20), .ZN(n_0_411));
   AOI222_X1 i_0_17_42 (.A1(n_0_390), .A2(n_0_378), .B1(n_0_391), .B2(n_0_346), 
      .C1(n_0_389), .C2(n_0_315), .ZN(n_0_17_21));
   INV_X1 i_0_17_43 (.A(n_0_17_21), .ZN(n_0_412));
   AOI222_X1 i_0_17_44 (.A1(n_0_390), .A2(n_0_379), .B1(n_0_391), .B2(n_0_347), 
      .C1(n_0_389), .C2(n_0_316), .ZN(n_0_17_22));
   INV_X1 i_0_17_45 (.A(n_0_17_22), .ZN(n_0_413));
   AOI222_X1 i_0_17_46 (.A1(n_0_390), .A2(n_0_380), .B1(n_0_391), .B2(n_0_348), 
      .C1(n_0_389), .C2(n_0_317), .ZN(n_0_17_23));
   INV_X1 i_0_17_47 (.A(n_0_17_23), .ZN(n_0_414));
   AOI222_X1 i_0_17_48 (.A1(n_0_390), .A2(n_0_381), .B1(n_0_391), .B2(n_0_349), 
      .C1(n_0_389), .C2(n_0_318), .ZN(n_0_17_24));
   INV_X1 i_0_17_49 (.A(n_0_17_24), .ZN(n_0_415));
   AOI222_X1 i_0_17_50 (.A1(n_0_390), .A2(n_0_382), .B1(n_0_391), .B2(n_0_350), 
      .C1(n_0_389), .C2(n_0_319), .ZN(n_0_17_25));
   INV_X1 i_0_17_51 (.A(n_0_17_25), .ZN(n_0_416));
   AOI222_X1 i_0_17_52 (.A1(n_0_390), .A2(n_0_383), .B1(n_0_391), .B2(n_0_351), 
      .C1(n_0_389), .C2(n_0_320), .ZN(n_0_17_26));
   INV_X1 i_0_17_53 (.A(n_0_17_26), .ZN(n_0_417));
   AOI222_X1 i_0_17_54 (.A1(n_0_390), .A2(n_0_384), .B1(n_0_391), .B2(n_0_352), 
      .C1(n_0_389), .C2(n_0_321), .ZN(n_0_17_27));
   INV_X1 i_0_17_55 (.A(n_0_17_27), .ZN(n_0_418));
   AOI222_X1 i_0_17_56 (.A1(n_0_390), .A2(n_0_385), .B1(n_0_391), .B2(n_0_353), 
      .C1(n_0_389), .C2(n_0_322), .ZN(n_0_17_28));
   INV_X1 i_0_17_57 (.A(n_0_17_28), .ZN(n_0_419));
   AOI222_X1 i_0_17_58 (.A1(n_0_390), .A2(n_0_386), .B1(n_0_391), .B2(n_0_354), 
      .C1(n_0_389), .C2(n_0_323), .ZN(n_0_17_29));
   INV_X1 i_0_17_59 (.A(n_0_17_29), .ZN(n_0_420));
   AND2_X1 i_0_17_60 (.A1(n_0_389), .A2(n_0_324), .ZN(n_0_17_30));
   AOI221_X1 i_0_17_61 (.A(n_0_17_30), .B1(n_0_390), .B2(n_0_387), .C1(n_0_391), 
      .C2(n_0_355), .ZN(n_0_17_31));
   INV_X1 i_0_17_62 (.A(n_0_17_31), .ZN(n_0_421));
   AOI221_X1 i_0_17_63 (.A(n_0_17_30), .B1(n_0_390), .B2(n_0_388), .C1(n_0_391), 
      .C2(n_0_356), .ZN(n_0_17_32));
   INV_X1 i_0_17_64 (.A(n_0_17_32), .ZN(n_0_422));
   datapath__0_16 i_0_18 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_9, 
      n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, n_0_415, 
      n_0_414, n_0_413, n_0_412, n_0_411, n_0_410, n_0_409, n_0_408, n_0_407, 
      n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, n_0_401, n_0_400, n_0_399, 
      n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, n_0_392}), .p_2({
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, n_0_444, n_0_443, n_0_442, n_0_441, n_0_440, n_0_439, 
      n_0_438, n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, n_0_432, n_0_431, 
      n_0_430, n_0_429, n_0_428, n_0_427, n_0_426, n_0_425, n_0_424, n_0_423}));
   datapath__0_17 i_0_19 (.multiplicand2(multiplicand2), .p_0({uc_10, n_0_422, 
      n_0_421, n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, n_0_415, n_0_414, 
      n_0_413, n_0_412, n_0_411, n_0_410, n_0_409, n_0_408, n_0_407, n_0_406, 
      n_0_405, n_0_404, n_0_403, n_0_402, n_0_401, n_0_400, n_0_399, n_0_398, 
      n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, n_0_392}), .p_1({n_0_486, 
      n_0_485, n_0_484, n_0_483, n_0_482, n_0_481, n_0_480, n_0_479, n_0_478, 
      n_0_477, n_0_476, n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, n_0_470, 
      n_0_469, n_0_468, n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, n_0_462, 
      n_0_461, n_0_460, n_0_459, n_0_458, n_0_457, n_0_456, n_0_455}));
   INV_X1 i_0_20_0 (.A(multiplier2[5]), .ZN(n_0_20_0));
   AND2_X1 i_0_20_1 (.A1(n_0_20_0), .A2(multiplier2[4]), .ZN(n_0_488));
   NOR2_X1 i_0_20_2 (.A1(n_0_20_0), .A2(multiplier2[4]), .ZN(n_0_489));
   NOR2_X1 i_0_20_3 (.A1(n_0_488), .A2(n_0_489), .ZN(n_0_487));
   AOI222_X1 i_0_21_0 (.A1(n_0_455), .A2(n_0_488), .B1(n_0_423), .B2(n_0_489), 
      .C1(n_0_392), .C2(n_0_487), .ZN(n_0_21_0));
   INV_X1 i_0_21_1 (.A(n_0_21_0), .ZN(product[5]));
   AOI222_X1 i_0_21_2 (.A1(n_0_488), .A2(n_0_456), .B1(n_0_489), .B2(n_0_424), 
      .C1(n_0_487), .C2(n_0_393), .ZN(n_0_21_1));
   INV_X1 i_0_21_3 (.A(n_0_21_1), .ZN(n_0_490));
   AOI222_X1 i_0_21_4 (.A1(n_0_488), .A2(n_0_457), .B1(n_0_489), .B2(n_0_425), 
      .C1(n_0_487), .C2(n_0_394), .ZN(n_0_21_2));
   INV_X1 i_0_21_5 (.A(n_0_21_2), .ZN(n_0_491));
   AOI222_X1 i_0_21_6 (.A1(n_0_488), .A2(n_0_458), .B1(n_0_489), .B2(n_0_426), 
      .C1(n_0_487), .C2(n_0_395), .ZN(n_0_21_3));
   INV_X1 i_0_21_7 (.A(n_0_21_3), .ZN(n_0_492));
   AOI222_X1 i_0_21_8 (.A1(n_0_488), .A2(n_0_459), .B1(n_0_489), .B2(n_0_427), 
      .C1(n_0_487), .C2(n_0_396), .ZN(n_0_21_4));
   INV_X1 i_0_21_9 (.A(n_0_21_4), .ZN(n_0_493));
   AOI222_X1 i_0_21_10 (.A1(n_0_488), .A2(n_0_460), .B1(n_0_489), .B2(n_0_428), 
      .C1(n_0_487), .C2(n_0_397), .ZN(n_0_21_5));
   INV_X1 i_0_21_11 (.A(n_0_21_5), .ZN(n_0_494));
   AOI222_X1 i_0_21_12 (.A1(n_0_488), .A2(n_0_461), .B1(n_0_489), .B2(n_0_429), 
      .C1(n_0_487), .C2(n_0_398), .ZN(n_0_21_6));
   INV_X1 i_0_21_13 (.A(n_0_21_6), .ZN(n_0_495));
   AOI222_X1 i_0_21_14 (.A1(n_0_488), .A2(n_0_462), .B1(n_0_489), .B2(n_0_430), 
      .C1(n_0_487), .C2(n_0_399), .ZN(n_0_21_7));
   INV_X1 i_0_21_15 (.A(n_0_21_7), .ZN(n_0_496));
   AOI222_X1 i_0_21_16 (.A1(n_0_488), .A2(n_0_463), .B1(n_0_489), .B2(n_0_431), 
      .C1(n_0_487), .C2(n_0_400), .ZN(n_0_21_8));
   INV_X1 i_0_21_17 (.A(n_0_21_8), .ZN(n_0_497));
   AOI222_X1 i_0_21_18 (.A1(n_0_488), .A2(n_0_464), .B1(n_0_489), .B2(n_0_432), 
      .C1(n_0_487), .C2(n_0_401), .ZN(n_0_21_9));
   INV_X1 i_0_21_19 (.A(n_0_21_9), .ZN(n_0_498));
   AOI222_X1 i_0_21_20 (.A1(n_0_488), .A2(n_0_465), .B1(n_0_489), .B2(n_0_433), 
      .C1(n_0_487), .C2(n_0_402), .ZN(n_0_21_10));
   INV_X1 i_0_21_21 (.A(n_0_21_10), .ZN(n_0_499));
   AOI222_X1 i_0_21_22 (.A1(n_0_488), .A2(n_0_466), .B1(n_0_489), .B2(n_0_434), 
      .C1(n_0_487), .C2(n_0_403), .ZN(n_0_21_11));
   INV_X1 i_0_21_23 (.A(n_0_21_11), .ZN(n_0_500));
   AOI222_X1 i_0_21_24 (.A1(n_0_488), .A2(n_0_467), .B1(n_0_489), .B2(n_0_435), 
      .C1(n_0_487), .C2(n_0_404), .ZN(n_0_21_12));
   INV_X1 i_0_21_25 (.A(n_0_21_12), .ZN(n_0_501));
   AOI222_X1 i_0_21_26 (.A1(n_0_488), .A2(n_0_468), .B1(n_0_489), .B2(n_0_436), 
      .C1(n_0_487), .C2(n_0_405), .ZN(n_0_21_13));
   INV_X1 i_0_21_27 (.A(n_0_21_13), .ZN(n_0_502));
   AOI222_X1 i_0_21_28 (.A1(n_0_488), .A2(n_0_469), .B1(n_0_489), .B2(n_0_437), 
      .C1(n_0_487), .C2(n_0_406), .ZN(n_0_21_14));
   INV_X1 i_0_21_29 (.A(n_0_21_14), .ZN(n_0_503));
   AOI222_X1 i_0_21_30 (.A1(n_0_488), .A2(n_0_470), .B1(n_0_489), .B2(n_0_438), 
      .C1(n_0_487), .C2(n_0_407), .ZN(n_0_21_15));
   INV_X1 i_0_21_31 (.A(n_0_21_15), .ZN(n_0_504));
   AOI222_X1 i_0_21_32 (.A1(n_0_488), .A2(n_0_471), .B1(n_0_489), .B2(n_0_439), 
      .C1(n_0_487), .C2(n_0_408), .ZN(n_0_21_16));
   INV_X1 i_0_21_33 (.A(n_0_21_16), .ZN(n_0_505));
   AOI222_X1 i_0_21_34 (.A1(n_0_488), .A2(n_0_472), .B1(n_0_489), .B2(n_0_440), 
      .C1(n_0_487), .C2(n_0_409), .ZN(n_0_21_17));
   INV_X1 i_0_21_35 (.A(n_0_21_17), .ZN(n_0_506));
   AOI222_X1 i_0_21_36 (.A1(n_0_488), .A2(n_0_473), .B1(n_0_489), .B2(n_0_441), 
      .C1(n_0_487), .C2(n_0_410), .ZN(n_0_21_18));
   INV_X1 i_0_21_37 (.A(n_0_21_18), .ZN(n_0_507));
   AOI222_X1 i_0_21_38 (.A1(n_0_488), .A2(n_0_474), .B1(n_0_489), .B2(n_0_442), 
      .C1(n_0_487), .C2(n_0_411), .ZN(n_0_21_19));
   INV_X1 i_0_21_39 (.A(n_0_21_19), .ZN(n_0_508));
   AOI222_X1 i_0_21_40 (.A1(n_0_488), .A2(n_0_475), .B1(n_0_489), .B2(n_0_443), 
      .C1(n_0_487), .C2(n_0_412), .ZN(n_0_21_20));
   INV_X1 i_0_21_41 (.A(n_0_21_20), .ZN(n_0_509));
   AOI222_X1 i_0_21_42 (.A1(n_0_488), .A2(n_0_476), .B1(n_0_489), .B2(n_0_444), 
      .C1(n_0_487), .C2(n_0_413), .ZN(n_0_21_21));
   INV_X1 i_0_21_43 (.A(n_0_21_21), .ZN(n_0_510));
   AOI222_X1 i_0_21_44 (.A1(n_0_488), .A2(n_0_477), .B1(n_0_489), .B2(n_0_445), 
      .C1(n_0_487), .C2(n_0_414), .ZN(n_0_21_22));
   INV_X1 i_0_21_45 (.A(n_0_21_22), .ZN(n_0_511));
   AOI222_X1 i_0_21_46 (.A1(n_0_488), .A2(n_0_478), .B1(n_0_489), .B2(n_0_446), 
      .C1(n_0_487), .C2(n_0_415), .ZN(n_0_21_23));
   INV_X1 i_0_21_47 (.A(n_0_21_23), .ZN(n_0_512));
   AOI222_X1 i_0_21_48 (.A1(n_0_488), .A2(n_0_479), .B1(n_0_489), .B2(n_0_447), 
      .C1(n_0_487), .C2(n_0_416), .ZN(n_0_21_24));
   INV_X1 i_0_21_49 (.A(n_0_21_24), .ZN(n_0_513));
   AOI222_X1 i_0_21_50 (.A1(n_0_488), .A2(n_0_480), .B1(n_0_489), .B2(n_0_448), 
      .C1(n_0_487), .C2(n_0_417), .ZN(n_0_21_25));
   INV_X1 i_0_21_51 (.A(n_0_21_25), .ZN(n_0_514));
   AOI222_X1 i_0_21_52 (.A1(n_0_488), .A2(n_0_481), .B1(n_0_489), .B2(n_0_449), 
      .C1(n_0_487), .C2(n_0_418), .ZN(n_0_21_26));
   INV_X1 i_0_21_53 (.A(n_0_21_26), .ZN(n_0_515));
   AOI222_X1 i_0_21_54 (.A1(n_0_488), .A2(n_0_482), .B1(n_0_489), .B2(n_0_450), 
      .C1(n_0_487), .C2(n_0_419), .ZN(n_0_21_27));
   INV_X1 i_0_21_55 (.A(n_0_21_27), .ZN(n_0_516));
   AOI222_X1 i_0_21_56 (.A1(n_0_488), .A2(n_0_483), .B1(n_0_489), .B2(n_0_451), 
      .C1(n_0_487), .C2(n_0_420), .ZN(n_0_21_28));
   INV_X1 i_0_21_57 (.A(n_0_21_28), .ZN(n_0_517));
   AOI222_X1 i_0_21_58 (.A1(n_0_488), .A2(n_0_484), .B1(n_0_489), .B2(n_0_452), 
      .C1(n_0_487), .C2(n_0_421), .ZN(n_0_21_29));
   INV_X1 i_0_21_59 (.A(n_0_21_29), .ZN(n_0_518));
   AND2_X1 i_0_21_60 (.A1(n_0_487), .A2(n_0_422), .ZN(n_0_21_30));
   AOI221_X1 i_0_21_61 (.A(n_0_21_30), .B1(n_0_488), .B2(n_0_485), .C1(n_0_489), 
      .C2(n_0_453), .ZN(n_0_21_31));
   INV_X1 i_0_21_62 (.A(n_0_21_31), .ZN(n_0_519));
   AOI221_X1 i_0_21_63 (.A(n_0_21_30), .B1(n_0_488), .B2(n_0_486), .C1(n_0_489), 
      .C2(n_0_454), .ZN(n_0_21_32));
   INV_X1 i_0_21_64 (.A(n_0_21_32), .ZN(n_0_520));
   datapath__0_20 i_0_22 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_11, 
      n_0_520, n_0_519, n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, 
      n_0_512, n_0_511, n_0_510, n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, 
      n_0_504, n_0_503, n_0_502, n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, 
      n_0_496, n_0_495, n_0_494, n_0_493, n_0_492, n_0_491, n_0_490}), .p_2({
      n_0_552, n_0_551, n_0_550, n_0_549, n_0_548, n_0_547, n_0_546, n_0_545, 
      n_0_544, n_0_543, n_0_542, n_0_541, n_0_540, n_0_539, n_0_538, n_0_537, 
      n_0_536, n_0_535, n_0_534, n_0_533, n_0_532, n_0_531, n_0_530, n_0_529, 
      n_0_528, n_0_527, n_0_526, n_0_525, n_0_524, n_0_523, n_0_522, n_0_521}));
   datapath__0_21 i_0_23 (.multiplicand2(multiplicand2), .p_0({uc_12, n_0_520, 
      n_0_519, n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, n_0_512, 
      n_0_511, n_0_510, n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, n_0_504, 
      n_0_503, n_0_502, n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, n_0_496, 
      n_0_495, n_0_494, n_0_493, n_0_492, n_0_491, n_0_490}), .p_1({n_0_584, 
      n_0_583, n_0_582, n_0_581, n_0_580, n_0_579, n_0_578, n_0_577, n_0_576, 
      n_0_575, n_0_574, n_0_573, n_0_572, n_0_571, n_0_570, n_0_569, n_0_568, 
      n_0_567, n_0_566, n_0_565, n_0_564, n_0_563, n_0_562, n_0_561, n_0_560, 
      n_0_559, n_0_558, n_0_557, n_0_556, n_0_555, n_0_554, n_0_553}));
   INV_X1 i_0_24_0 (.A(multiplier2[6]), .ZN(n_0_24_0));
   AND2_X1 i_0_24_1 (.A1(n_0_24_0), .A2(multiplier2[5]), .ZN(n_0_586));
   NOR2_X1 i_0_24_2 (.A1(n_0_24_0), .A2(multiplier2[5]), .ZN(n_0_587));
   NOR2_X1 i_0_24_3 (.A1(n_0_586), .A2(n_0_587), .ZN(n_0_585));
   AOI222_X1 i_0_25_0 (.A1(n_0_553), .A2(n_0_586), .B1(n_0_521), .B2(n_0_587), 
      .C1(n_0_490), .C2(n_0_585), .ZN(n_0_25_0));
   INV_X1 i_0_25_1 (.A(n_0_25_0), .ZN(product[6]));
   AOI222_X1 i_0_25_2 (.A1(n_0_586), .A2(n_0_554), .B1(n_0_587), .B2(n_0_522), 
      .C1(n_0_585), .C2(n_0_491), .ZN(n_0_25_1));
   INV_X1 i_0_25_3 (.A(n_0_25_1), .ZN(n_0_588));
   AOI222_X1 i_0_25_4 (.A1(n_0_586), .A2(n_0_555), .B1(n_0_587), .B2(n_0_523), 
      .C1(n_0_585), .C2(n_0_492), .ZN(n_0_25_2));
   INV_X1 i_0_25_5 (.A(n_0_25_2), .ZN(n_0_589));
   AOI222_X1 i_0_25_6 (.A1(n_0_586), .A2(n_0_556), .B1(n_0_587), .B2(n_0_524), 
      .C1(n_0_585), .C2(n_0_493), .ZN(n_0_25_3));
   INV_X1 i_0_25_7 (.A(n_0_25_3), .ZN(n_0_590));
   AOI222_X1 i_0_25_8 (.A1(n_0_586), .A2(n_0_557), .B1(n_0_587), .B2(n_0_525), 
      .C1(n_0_585), .C2(n_0_494), .ZN(n_0_25_4));
   INV_X1 i_0_25_9 (.A(n_0_25_4), .ZN(n_0_591));
   AOI222_X1 i_0_25_10 (.A1(n_0_586), .A2(n_0_558), .B1(n_0_587), .B2(n_0_526), 
      .C1(n_0_585), .C2(n_0_495), .ZN(n_0_25_5));
   INV_X1 i_0_25_11 (.A(n_0_25_5), .ZN(n_0_592));
   AOI222_X1 i_0_25_12 (.A1(n_0_586), .A2(n_0_559), .B1(n_0_587), .B2(n_0_527), 
      .C1(n_0_585), .C2(n_0_496), .ZN(n_0_25_6));
   INV_X1 i_0_25_13 (.A(n_0_25_6), .ZN(n_0_593));
   AOI222_X1 i_0_25_14 (.A1(n_0_586), .A2(n_0_560), .B1(n_0_587), .B2(n_0_528), 
      .C1(n_0_585), .C2(n_0_497), .ZN(n_0_25_7));
   INV_X1 i_0_25_15 (.A(n_0_25_7), .ZN(n_0_594));
   AOI222_X1 i_0_25_16 (.A1(n_0_586), .A2(n_0_561), .B1(n_0_587), .B2(n_0_529), 
      .C1(n_0_585), .C2(n_0_498), .ZN(n_0_25_8));
   INV_X1 i_0_25_17 (.A(n_0_25_8), .ZN(n_0_595));
   AOI222_X1 i_0_25_18 (.A1(n_0_586), .A2(n_0_562), .B1(n_0_587), .B2(n_0_530), 
      .C1(n_0_585), .C2(n_0_499), .ZN(n_0_25_9));
   INV_X1 i_0_25_19 (.A(n_0_25_9), .ZN(n_0_596));
   AOI222_X1 i_0_25_20 (.A1(n_0_586), .A2(n_0_563), .B1(n_0_587), .B2(n_0_531), 
      .C1(n_0_585), .C2(n_0_500), .ZN(n_0_25_10));
   INV_X1 i_0_25_21 (.A(n_0_25_10), .ZN(n_0_597));
   AOI222_X1 i_0_25_22 (.A1(n_0_586), .A2(n_0_564), .B1(n_0_587), .B2(n_0_532), 
      .C1(n_0_585), .C2(n_0_501), .ZN(n_0_25_11));
   INV_X1 i_0_25_23 (.A(n_0_25_11), .ZN(n_0_598));
   AOI222_X1 i_0_25_24 (.A1(n_0_586), .A2(n_0_565), .B1(n_0_587), .B2(n_0_533), 
      .C1(n_0_585), .C2(n_0_502), .ZN(n_0_25_12));
   INV_X1 i_0_25_25 (.A(n_0_25_12), .ZN(n_0_599));
   AOI222_X1 i_0_25_26 (.A1(n_0_586), .A2(n_0_566), .B1(n_0_587), .B2(n_0_534), 
      .C1(n_0_585), .C2(n_0_503), .ZN(n_0_25_13));
   INV_X1 i_0_25_27 (.A(n_0_25_13), .ZN(n_0_600));
   AOI222_X1 i_0_25_28 (.A1(n_0_586), .A2(n_0_567), .B1(n_0_587), .B2(n_0_535), 
      .C1(n_0_585), .C2(n_0_504), .ZN(n_0_25_14));
   INV_X1 i_0_25_29 (.A(n_0_25_14), .ZN(n_0_601));
   AOI222_X1 i_0_25_30 (.A1(n_0_586), .A2(n_0_568), .B1(n_0_587), .B2(n_0_536), 
      .C1(n_0_585), .C2(n_0_505), .ZN(n_0_25_15));
   INV_X1 i_0_25_31 (.A(n_0_25_15), .ZN(n_0_602));
   AOI222_X1 i_0_25_32 (.A1(n_0_586), .A2(n_0_569), .B1(n_0_587), .B2(n_0_537), 
      .C1(n_0_585), .C2(n_0_506), .ZN(n_0_25_16));
   INV_X1 i_0_25_33 (.A(n_0_25_16), .ZN(n_0_603));
   AOI222_X1 i_0_25_34 (.A1(n_0_586), .A2(n_0_570), .B1(n_0_587), .B2(n_0_538), 
      .C1(n_0_585), .C2(n_0_507), .ZN(n_0_25_17));
   INV_X1 i_0_25_35 (.A(n_0_25_17), .ZN(n_0_604));
   AOI222_X1 i_0_25_36 (.A1(n_0_586), .A2(n_0_571), .B1(n_0_587), .B2(n_0_539), 
      .C1(n_0_585), .C2(n_0_508), .ZN(n_0_25_18));
   INV_X1 i_0_25_37 (.A(n_0_25_18), .ZN(n_0_605));
   AOI222_X1 i_0_25_38 (.A1(n_0_586), .A2(n_0_572), .B1(n_0_587), .B2(n_0_540), 
      .C1(n_0_585), .C2(n_0_509), .ZN(n_0_25_19));
   INV_X1 i_0_25_39 (.A(n_0_25_19), .ZN(n_0_606));
   AOI222_X1 i_0_25_40 (.A1(n_0_586), .A2(n_0_573), .B1(n_0_587), .B2(n_0_541), 
      .C1(n_0_585), .C2(n_0_510), .ZN(n_0_25_20));
   INV_X1 i_0_25_41 (.A(n_0_25_20), .ZN(n_0_607));
   AOI222_X1 i_0_25_42 (.A1(n_0_586), .A2(n_0_574), .B1(n_0_587), .B2(n_0_542), 
      .C1(n_0_585), .C2(n_0_511), .ZN(n_0_25_21));
   INV_X1 i_0_25_43 (.A(n_0_25_21), .ZN(n_0_608));
   AOI222_X1 i_0_25_44 (.A1(n_0_586), .A2(n_0_575), .B1(n_0_587), .B2(n_0_543), 
      .C1(n_0_585), .C2(n_0_512), .ZN(n_0_25_22));
   INV_X1 i_0_25_45 (.A(n_0_25_22), .ZN(n_0_609));
   AOI222_X1 i_0_25_46 (.A1(n_0_586), .A2(n_0_576), .B1(n_0_587), .B2(n_0_544), 
      .C1(n_0_585), .C2(n_0_513), .ZN(n_0_25_23));
   INV_X1 i_0_25_47 (.A(n_0_25_23), .ZN(n_0_610));
   AOI222_X1 i_0_25_48 (.A1(n_0_586), .A2(n_0_577), .B1(n_0_587), .B2(n_0_545), 
      .C1(n_0_585), .C2(n_0_514), .ZN(n_0_25_24));
   INV_X1 i_0_25_49 (.A(n_0_25_24), .ZN(n_0_611));
   AOI222_X1 i_0_25_50 (.A1(n_0_586), .A2(n_0_578), .B1(n_0_587), .B2(n_0_546), 
      .C1(n_0_585), .C2(n_0_515), .ZN(n_0_25_25));
   INV_X1 i_0_25_51 (.A(n_0_25_25), .ZN(n_0_612));
   AOI222_X1 i_0_25_52 (.A1(n_0_586), .A2(n_0_579), .B1(n_0_587), .B2(n_0_547), 
      .C1(n_0_585), .C2(n_0_516), .ZN(n_0_25_26));
   INV_X1 i_0_25_53 (.A(n_0_25_26), .ZN(n_0_613));
   AOI222_X1 i_0_25_54 (.A1(n_0_586), .A2(n_0_580), .B1(n_0_587), .B2(n_0_548), 
      .C1(n_0_585), .C2(n_0_517), .ZN(n_0_25_27));
   INV_X1 i_0_25_55 (.A(n_0_25_27), .ZN(n_0_614));
   AOI222_X1 i_0_25_56 (.A1(n_0_586), .A2(n_0_581), .B1(n_0_587), .B2(n_0_549), 
      .C1(n_0_585), .C2(n_0_518), .ZN(n_0_25_28));
   INV_X1 i_0_25_57 (.A(n_0_25_28), .ZN(n_0_615));
   AOI222_X1 i_0_25_58 (.A1(n_0_586), .A2(n_0_582), .B1(n_0_587), .B2(n_0_550), 
      .C1(n_0_585), .C2(n_0_519), .ZN(n_0_25_29));
   INV_X1 i_0_25_59 (.A(n_0_25_29), .ZN(n_0_616));
   AND2_X1 i_0_25_60 (.A1(n_0_585), .A2(n_0_520), .ZN(n_0_25_30));
   AOI221_X1 i_0_25_61 (.A(n_0_25_30), .B1(n_0_586), .B2(n_0_583), .C1(n_0_587), 
      .C2(n_0_551), .ZN(n_0_25_31));
   INV_X1 i_0_25_62 (.A(n_0_25_31), .ZN(n_0_617));
   AOI221_X1 i_0_25_63 (.A(n_0_25_30), .B1(n_0_586), .B2(n_0_584), .C1(n_0_587), 
      .C2(n_0_552), .ZN(n_0_25_32));
   INV_X1 i_0_25_64 (.A(n_0_25_32), .ZN(n_0_618));
   datapath__0_24 i_0_26 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_13, 
      n_0_618, n_0_617, n_0_616, n_0_615, n_0_614, n_0_613, n_0_612, n_0_611, 
      n_0_610, n_0_609, n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, n_0_603, 
      n_0_602, n_0_601, n_0_600, n_0_599, n_0_598, n_0_597, n_0_596, n_0_595, 
      n_0_594, n_0_593, n_0_592, n_0_591, n_0_590, n_0_589, n_0_588}), .p_2({
      n_0_650, n_0_649, n_0_648, n_0_647, n_0_646, n_0_645, n_0_644, n_0_643, 
      n_0_642, n_0_641, n_0_640, n_0_639, n_0_638, n_0_637, n_0_636, n_0_635, 
      n_0_634, n_0_633, n_0_632, n_0_631, n_0_630, n_0_629, n_0_628, n_0_627, 
      n_0_626, n_0_625, n_0_624, n_0_623, n_0_622, n_0_621, n_0_620, n_0_619}));
   datapath__0_25 i_0_27 (.multiplicand2(multiplicand2), .p_0({uc_14, n_0_618, 
      n_0_617, n_0_616, n_0_615, n_0_614, n_0_613, n_0_612, n_0_611, n_0_610, 
      n_0_609, n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, n_0_603, n_0_602, 
      n_0_601, n_0_600, n_0_599, n_0_598, n_0_597, n_0_596, n_0_595, n_0_594, 
      n_0_593, n_0_592, n_0_591, n_0_590, n_0_589, n_0_588}), .p_1({n_0_682, 
      n_0_681, n_0_680, n_0_679, n_0_678, n_0_677, n_0_676, n_0_675, n_0_674, 
      n_0_673, n_0_672, n_0_671, n_0_670, n_0_669, n_0_668, n_0_667, n_0_666, 
      n_0_665, n_0_664, n_0_663, n_0_662, n_0_661, n_0_660, n_0_659, n_0_658, 
      n_0_657, n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, n_0_651}));
   INV_X1 i_0_28_0 (.A(multiplier2[7]), .ZN(n_0_28_0));
   AND2_X1 i_0_28_1 (.A1(n_0_28_0), .A2(multiplier2[6]), .ZN(n_0_684));
   NOR2_X1 i_0_28_2 (.A1(n_0_28_0), .A2(multiplier2[6]), .ZN(n_0_685));
   NOR2_X1 i_0_28_3 (.A1(n_0_684), .A2(n_0_685), .ZN(n_0_683));
   AOI222_X1 i_0_29_0 (.A1(n_0_651), .A2(n_0_684), .B1(n_0_619), .B2(n_0_685), 
      .C1(n_0_588), .C2(n_0_683), .ZN(n_0_29_0));
   INV_X1 i_0_29_1 (.A(n_0_29_0), .ZN(product[7]));
   AOI222_X1 i_0_29_2 (.A1(n_0_684), .A2(n_0_652), .B1(n_0_685), .B2(n_0_620), 
      .C1(n_0_683), .C2(n_0_589), .ZN(n_0_29_1));
   INV_X1 i_0_29_3 (.A(n_0_29_1), .ZN(n_0_686));
   AOI222_X1 i_0_29_4 (.A1(n_0_684), .A2(n_0_653), .B1(n_0_685), .B2(n_0_621), 
      .C1(n_0_683), .C2(n_0_590), .ZN(n_0_29_2));
   INV_X1 i_0_29_5 (.A(n_0_29_2), .ZN(n_0_687));
   AOI222_X1 i_0_29_6 (.A1(n_0_684), .A2(n_0_654), .B1(n_0_685), .B2(n_0_622), 
      .C1(n_0_683), .C2(n_0_591), .ZN(n_0_29_3));
   INV_X1 i_0_29_7 (.A(n_0_29_3), .ZN(n_0_688));
   AOI222_X1 i_0_29_8 (.A1(n_0_684), .A2(n_0_655), .B1(n_0_685), .B2(n_0_623), 
      .C1(n_0_683), .C2(n_0_592), .ZN(n_0_29_4));
   INV_X1 i_0_29_9 (.A(n_0_29_4), .ZN(n_0_689));
   AOI222_X1 i_0_29_10 (.A1(n_0_684), .A2(n_0_656), .B1(n_0_685), .B2(n_0_624), 
      .C1(n_0_683), .C2(n_0_593), .ZN(n_0_29_5));
   INV_X1 i_0_29_11 (.A(n_0_29_5), .ZN(n_0_690));
   AOI222_X1 i_0_29_12 (.A1(n_0_684), .A2(n_0_657), .B1(n_0_685), .B2(n_0_625), 
      .C1(n_0_683), .C2(n_0_594), .ZN(n_0_29_6));
   INV_X1 i_0_29_13 (.A(n_0_29_6), .ZN(n_0_691));
   AOI222_X1 i_0_29_14 (.A1(n_0_684), .A2(n_0_658), .B1(n_0_685), .B2(n_0_626), 
      .C1(n_0_683), .C2(n_0_595), .ZN(n_0_29_7));
   INV_X1 i_0_29_15 (.A(n_0_29_7), .ZN(n_0_692));
   AOI222_X1 i_0_29_16 (.A1(n_0_684), .A2(n_0_659), .B1(n_0_685), .B2(n_0_627), 
      .C1(n_0_683), .C2(n_0_596), .ZN(n_0_29_8));
   INV_X1 i_0_29_17 (.A(n_0_29_8), .ZN(n_0_693));
   AOI222_X1 i_0_29_18 (.A1(n_0_684), .A2(n_0_660), .B1(n_0_685), .B2(n_0_628), 
      .C1(n_0_683), .C2(n_0_597), .ZN(n_0_29_9));
   INV_X1 i_0_29_19 (.A(n_0_29_9), .ZN(n_0_694));
   AOI222_X1 i_0_29_20 (.A1(n_0_684), .A2(n_0_661), .B1(n_0_685), .B2(n_0_629), 
      .C1(n_0_683), .C2(n_0_598), .ZN(n_0_29_10));
   INV_X1 i_0_29_21 (.A(n_0_29_10), .ZN(n_0_695));
   AOI222_X1 i_0_29_22 (.A1(n_0_684), .A2(n_0_662), .B1(n_0_685), .B2(n_0_630), 
      .C1(n_0_683), .C2(n_0_599), .ZN(n_0_29_11));
   INV_X1 i_0_29_23 (.A(n_0_29_11), .ZN(n_0_696));
   AOI222_X1 i_0_29_24 (.A1(n_0_684), .A2(n_0_663), .B1(n_0_685), .B2(n_0_631), 
      .C1(n_0_683), .C2(n_0_600), .ZN(n_0_29_12));
   INV_X1 i_0_29_25 (.A(n_0_29_12), .ZN(n_0_697));
   AOI222_X1 i_0_29_26 (.A1(n_0_684), .A2(n_0_664), .B1(n_0_685), .B2(n_0_632), 
      .C1(n_0_683), .C2(n_0_601), .ZN(n_0_29_13));
   INV_X1 i_0_29_27 (.A(n_0_29_13), .ZN(n_0_698));
   AOI222_X1 i_0_29_28 (.A1(n_0_684), .A2(n_0_665), .B1(n_0_685), .B2(n_0_633), 
      .C1(n_0_683), .C2(n_0_602), .ZN(n_0_29_14));
   INV_X1 i_0_29_29 (.A(n_0_29_14), .ZN(n_0_699));
   AOI222_X1 i_0_29_30 (.A1(n_0_684), .A2(n_0_666), .B1(n_0_685), .B2(n_0_634), 
      .C1(n_0_683), .C2(n_0_603), .ZN(n_0_29_15));
   INV_X1 i_0_29_31 (.A(n_0_29_15), .ZN(n_0_700));
   AOI222_X1 i_0_29_32 (.A1(n_0_684), .A2(n_0_667), .B1(n_0_685), .B2(n_0_635), 
      .C1(n_0_683), .C2(n_0_604), .ZN(n_0_29_16));
   INV_X1 i_0_29_33 (.A(n_0_29_16), .ZN(n_0_701));
   AOI222_X1 i_0_29_34 (.A1(n_0_684), .A2(n_0_668), .B1(n_0_685), .B2(n_0_636), 
      .C1(n_0_683), .C2(n_0_605), .ZN(n_0_29_17));
   INV_X1 i_0_29_35 (.A(n_0_29_17), .ZN(n_0_702));
   AOI222_X1 i_0_29_36 (.A1(n_0_684), .A2(n_0_669), .B1(n_0_685), .B2(n_0_637), 
      .C1(n_0_683), .C2(n_0_606), .ZN(n_0_29_18));
   INV_X1 i_0_29_37 (.A(n_0_29_18), .ZN(n_0_703));
   AOI222_X1 i_0_29_38 (.A1(n_0_684), .A2(n_0_670), .B1(n_0_685), .B2(n_0_638), 
      .C1(n_0_683), .C2(n_0_607), .ZN(n_0_29_19));
   INV_X1 i_0_29_39 (.A(n_0_29_19), .ZN(n_0_704));
   AOI222_X1 i_0_29_40 (.A1(n_0_684), .A2(n_0_671), .B1(n_0_685), .B2(n_0_639), 
      .C1(n_0_683), .C2(n_0_608), .ZN(n_0_29_20));
   INV_X1 i_0_29_41 (.A(n_0_29_20), .ZN(n_0_705));
   AOI222_X1 i_0_29_42 (.A1(n_0_684), .A2(n_0_672), .B1(n_0_685), .B2(n_0_640), 
      .C1(n_0_683), .C2(n_0_609), .ZN(n_0_29_21));
   INV_X1 i_0_29_43 (.A(n_0_29_21), .ZN(n_0_706));
   AOI222_X1 i_0_29_44 (.A1(n_0_684), .A2(n_0_673), .B1(n_0_685), .B2(n_0_641), 
      .C1(n_0_683), .C2(n_0_610), .ZN(n_0_29_22));
   INV_X1 i_0_29_45 (.A(n_0_29_22), .ZN(n_0_707));
   AOI222_X1 i_0_29_46 (.A1(n_0_684), .A2(n_0_674), .B1(n_0_685), .B2(n_0_642), 
      .C1(n_0_683), .C2(n_0_611), .ZN(n_0_29_23));
   INV_X1 i_0_29_47 (.A(n_0_29_23), .ZN(n_0_708));
   AOI222_X1 i_0_29_48 (.A1(n_0_684), .A2(n_0_675), .B1(n_0_685), .B2(n_0_643), 
      .C1(n_0_683), .C2(n_0_612), .ZN(n_0_29_24));
   INV_X1 i_0_29_49 (.A(n_0_29_24), .ZN(n_0_709));
   AOI222_X1 i_0_29_50 (.A1(n_0_684), .A2(n_0_676), .B1(n_0_685), .B2(n_0_644), 
      .C1(n_0_683), .C2(n_0_613), .ZN(n_0_29_25));
   INV_X1 i_0_29_51 (.A(n_0_29_25), .ZN(n_0_710));
   AOI222_X1 i_0_29_52 (.A1(n_0_684), .A2(n_0_677), .B1(n_0_685), .B2(n_0_645), 
      .C1(n_0_683), .C2(n_0_614), .ZN(n_0_29_26));
   INV_X1 i_0_29_53 (.A(n_0_29_26), .ZN(n_0_711));
   AOI222_X1 i_0_29_54 (.A1(n_0_684), .A2(n_0_678), .B1(n_0_685), .B2(n_0_646), 
      .C1(n_0_683), .C2(n_0_615), .ZN(n_0_29_27));
   INV_X1 i_0_29_55 (.A(n_0_29_27), .ZN(n_0_712));
   AOI222_X1 i_0_29_56 (.A1(n_0_684), .A2(n_0_679), .B1(n_0_685), .B2(n_0_647), 
      .C1(n_0_683), .C2(n_0_616), .ZN(n_0_29_28));
   INV_X1 i_0_29_57 (.A(n_0_29_28), .ZN(n_0_713));
   AOI222_X1 i_0_29_58 (.A1(n_0_684), .A2(n_0_680), .B1(n_0_685), .B2(n_0_648), 
      .C1(n_0_683), .C2(n_0_617), .ZN(n_0_29_29));
   INV_X1 i_0_29_59 (.A(n_0_29_29), .ZN(n_0_714));
   AND2_X1 i_0_29_60 (.A1(n_0_683), .A2(n_0_618), .ZN(n_0_29_30));
   AOI221_X1 i_0_29_61 (.A(n_0_29_30), .B1(n_0_684), .B2(n_0_681), .C1(n_0_685), 
      .C2(n_0_649), .ZN(n_0_29_31));
   INV_X1 i_0_29_62 (.A(n_0_29_31), .ZN(n_0_715));
   AOI221_X1 i_0_29_63 (.A(n_0_29_30), .B1(n_0_684), .B2(n_0_682), .C1(n_0_685), 
      .C2(n_0_650), .ZN(n_0_29_32));
   INV_X1 i_0_29_64 (.A(n_0_29_32), .ZN(n_0_716));
   datapath__0_28 i_0_30 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_15, 
      n_0_716, n_0_715, n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, 
      n_0_708, n_0_707, n_0_706, n_0_705, n_0_704, n_0_703, n_0_702, n_0_701, 
      n_0_700, n_0_699, n_0_698, n_0_697, n_0_696, n_0_695, n_0_694, n_0_693, 
      n_0_692, n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686}), .p_2({
      n_0_748, n_0_747, n_0_746, n_0_745, n_0_744, n_0_743, n_0_742, n_0_741, 
      n_0_740, n_0_739, n_0_738, n_0_737, n_0_736, n_0_735, n_0_734, n_0_733, 
      n_0_732, n_0_731, n_0_730, n_0_729, n_0_728, n_0_727, n_0_726, n_0_725, 
      n_0_724, n_0_723, n_0_722, n_0_721, n_0_720, n_0_719, n_0_718, n_0_717}));
   datapath__0_29 i_0_31 (.multiplicand2(multiplicand2), .p_0({uc_16, n_0_716, 
      n_0_715, n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, 
      n_0_707, n_0_706, n_0_705, n_0_704, n_0_703, n_0_702, n_0_701, n_0_700, 
      n_0_699, n_0_698, n_0_697, n_0_696, n_0_695, n_0_694, n_0_693, n_0_692, 
      n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686}), .p_1({n_0_780, 
      n_0_779, n_0_778, n_0_777, n_0_776, n_0_775, n_0_774, n_0_773, n_0_772, 
      n_0_771, n_0_770, n_0_769, n_0_768, n_0_767, n_0_766, n_0_765, n_0_764, 
      n_0_763, n_0_762, n_0_761, n_0_760, n_0_759, n_0_758, n_0_757, n_0_756, 
      n_0_755, n_0_754, n_0_753, n_0_752, n_0_751, n_0_750, n_0_749}));
   INV_X1 i_0_32_0 (.A(multiplier2[8]), .ZN(n_0_32_0));
   AND2_X1 i_0_32_1 (.A1(n_0_32_0), .A2(multiplier2[7]), .ZN(n_0_782));
   NOR2_X1 i_0_32_2 (.A1(n_0_32_0), .A2(multiplier2[7]), .ZN(n_0_783));
   NOR2_X1 i_0_32_3 (.A1(n_0_782), .A2(n_0_783), .ZN(n_0_781));
   AOI222_X1 i_0_33_0 (.A1(n_0_749), .A2(n_0_782), .B1(n_0_717), .B2(n_0_783), 
      .C1(n_0_686), .C2(n_0_781), .ZN(n_0_33_0));
   INV_X1 i_0_33_1 (.A(n_0_33_0), .ZN(product[8]));
   AOI222_X1 i_0_33_2 (.A1(n_0_782), .A2(n_0_750), .B1(n_0_783), .B2(n_0_718), 
      .C1(n_0_781), .C2(n_0_687), .ZN(n_0_33_1));
   INV_X1 i_0_33_3 (.A(n_0_33_1), .ZN(n_0_784));
   AOI222_X1 i_0_33_4 (.A1(n_0_782), .A2(n_0_751), .B1(n_0_783), .B2(n_0_719), 
      .C1(n_0_781), .C2(n_0_688), .ZN(n_0_33_2));
   INV_X1 i_0_33_5 (.A(n_0_33_2), .ZN(n_0_785));
   AOI222_X1 i_0_33_6 (.A1(n_0_782), .A2(n_0_752), .B1(n_0_783), .B2(n_0_720), 
      .C1(n_0_781), .C2(n_0_689), .ZN(n_0_33_3));
   INV_X1 i_0_33_7 (.A(n_0_33_3), .ZN(n_0_786));
   AOI222_X1 i_0_33_8 (.A1(n_0_782), .A2(n_0_753), .B1(n_0_783), .B2(n_0_721), 
      .C1(n_0_781), .C2(n_0_690), .ZN(n_0_33_4));
   INV_X1 i_0_33_9 (.A(n_0_33_4), .ZN(n_0_787));
   AOI222_X1 i_0_33_10 (.A1(n_0_782), .A2(n_0_754), .B1(n_0_783), .B2(n_0_722), 
      .C1(n_0_781), .C2(n_0_691), .ZN(n_0_33_5));
   INV_X1 i_0_33_11 (.A(n_0_33_5), .ZN(n_0_788));
   AOI222_X1 i_0_33_12 (.A1(n_0_782), .A2(n_0_755), .B1(n_0_783), .B2(n_0_723), 
      .C1(n_0_781), .C2(n_0_692), .ZN(n_0_33_6));
   INV_X1 i_0_33_13 (.A(n_0_33_6), .ZN(n_0_789));
   AOI222_X1 i_0_33_14 (.A1(n_0_782), .A2(n_0_756), .B1(n_0_783), .B2(n_0_724), 
      .C1(n_0_781), .C2(n_0_693), .ZN(n_0_33_7));
   INV_X1 i_0_33_15 (.A(n_0_33_7), .ZN(n_0_790));
   AOI222_X1 i_0_33_16 (.A1(n_0_782), .A2(n_0_757), .B1(n_0_783), .B2(n_0_725), 
      .C1(n_0_781), .C2(n_0_694), .ZN(n_0_33_8));
   INV_X1 i_0_33_17 (.A(n_0_33_8), .ZN(n_0_791));
   AOI222_X1 i_0_33_18 (.A1(n_0_782), .A2(n_0_758), .B1(n_0_783), .B2(n_0_726), 
      .C1(n_0_781), .C2(n_0_695), .ZN(n_0_33_9));
   INV_X1 i_0_33_19 (.A(n_0_33_9), .ZN(n_0_792));
   AOI222_X1 i_0_33_20 (.A1(n_0_782), .A2(n_0_759), .B1(n_0_783), .B2(n_0_727), 
      .C1(n_0_781), .C2(n_0_696), .ZN(n_0_33_10));
   INV_X1 i_0_33_21 (.A(n_0_33_10), .ZN(n_0_793));
   AOI222_X1 i_0_33_22 (.A1(n_0_782), .A2(n_0_760), .B1(n_0_783), .B2(n_0_728), 
      .C1(n_0_781), .C2(n_0_697), .ZN(n_0_33_11));
   INV_X1 i_0_33_23 (.A(n_0_33_11), .ZN(n_0_794));
   AOI222_X1 i_0_33_24 (.A1(n_0_782), .A2(n_0_761), .B1(n_0_783), .B2(n_0_729), 
      .C1(n_0_781), .C2(n_0_698), .ZN(n_0_33_12));
   INV_X1 i_0_33_25 (.A(n_0_33_12), .ZN(n_0_795));
   AOI222_X1 i_0_33_26 (.A1(n_0_782), .A2(n_0_762), .B1(n_0_783), .B2(n_0_730), 
      .C1(n_0_781), .C2(n_0_699), .ZN(n_0_33_13));
   INV_X1 i_0_33_27 (.A(n_0_33_13), .ZN(n_0_796));
   AOI222_X1 i_0_33_28 (.A1(n_0_782), .A2(n_0_763), .B1(n_0_783), .B2(n_0_731), 
      .C1(n_0_781), .C2(n_0_700), .ZN(n_0_33_14));
   INV_X1 i_0_33_29 (.A(n_0_33_14), .ZN(n_0_797));
   AOI222_X1 i_0_33_30 (.A1(n_0_782), .A2(n_0_764), .B1(n_0_783), .B2(n_0_732), 
      .C1(n_0_781), .C2(n_0_701), .ZN(n_0_33_15));
   INV_X1 i_0_33_31 (.A(n_0_33_15), .ZN(n_0_798));
   AOI222_X1 i_0_33_32 (.A1(n_0_782), .A2(n_0_765), .B1(n_0_783), .B2(n_0_733), 
      .C1(n_0_781), .C2(n_0_702), .ZN(n_0_33_16));
   INV_X1 i_0_33_33 (.A(n_0_33_16), .ZN(n_0_799));
   AOI222_X1 i_0_33_34 (.A1(n_0_782), .A2(n_0_766), .B1(n_0_783), .B2(n_0_734), 
      .C1(n_0_781), .C2(n_0_703), .ZN(n_0_33_17));
   INV_X1 i_0_33_35 (.A(n_0_33_17), .ZN(n_0_800));
   AOI222_X1 i_0_33_36 (.A1(n_0_782), .A2(n_0_767), .B1(n_0_783), .B2(n_0_735), 
      .C1(n_0_781), .C2(n_0_704), .ZN(n_0_33_18));
   INV_X1 i_0_33_37 (.A(n_0_33_18), .ZN(n_0_801));
   AOI222_X1 i_0_33_38 (.A1(n_0_782), .A2(n_0_768), .B1(n_0_783), .B2(n_0_736), 
      .C1(n_0_781), .C2(n_0_705), .ZN(n_0_33_19));
   INV_X1 i_0_33_39 (.A(n_0_33_19), .ZN(n_0_802));
   AOI222_X1 i_0_33_40 (.A1(n_0_782), .A2(n_0_769), .B1(n_0_783), .B2(n_0_737), 
      .C1(n_0_781), .C2(n_0_706), .ZN(n_0_33_20));
   INV_X1 i_0_33_41 (.A(n_0_33_20), .ZN(n_0_803));
   AOI222_X1 i_0_33_42 (.A1(n_0_782), .A2(n_0_770), .B1(n_0_783), .B2(n_0_738), 
      .C1(n_0_781), .C2(n_0_707), .ZN(n_0_33_21));
   INV_X1 i_0_33_43 (.A(n_0_33_21), .ZN(n_0_804));
   AOI222_X1 i_0_33_44 (.A1(n_0_782), .A2(n_0_771), .B1(n_0_783), .B2(n_0_739), 
      .C1(n_0_781), .C2(n_0_708), .ZN(n_0_33_22));
   INV_X1 i_0_33_45 (.A(n_0_33_22), .ZN(n_0_805));
   AOI222_X1 i_0_33_46 (.A1(n_0_782), .A2(n_0_772), .B1(n_0_783), .B2(n_0_740), 
      .C1(n_0_781), .C2(n_0_709), .ZN(n_0_33_23));
   INV_X1 i_0_33_47 (.A(n_0_33_23), .ZN(n_0_806));
   AOI222_X1 i_0_33_48 (.A1(n_0_782), .A2(n_0_773), .B1(n_0_783), .B2(n_0_741), 
      .C1(n_0_781), .C2(n_0_710), .ZN(n_0_33_24));
   INV_X1 i_0_33_49 (.A(n_0_33_24), .ZN(n_0_807));
   AOI222_X1 i_0_33_50 (.A1(n_0_782), .A2(n_0_774), .B1(n_0_783), .B2(n_0_742), 
      .C1(n_0_781), .C2(n_0_711), .ZN(n_0_33_25));
   INV_X1 i_0_33_51 (.A(n_0_33_25), .ZN(n_0_808));
   AOI222_X1 i_0_33_52 (.A1(n_0_782), .A2(n_0_775), .B1(n_0_783), .B2(n_0_743), 
      .C1(n_0_781), .C2(n_0_712), .ZN(n_0_33_26));
   INV_X1 i_0_33_53 (.A(n_0_33_26), .ZN(n_0_809));
   AOI222_X1 i_0_33_54 (.A1(n_0_782), .A2(n_0_776), .B1(n_0_783), .B2(n_0_744), 
      .C1(n_0_781), .C2(n_0_713), .ZN(n_0_33_27));
   INV_X1 i_0_33_55 (.A(n_0_33_27), .ZN(n_0_810));
   AOI222_X1 i_0_33_56 (.A1(n_0_782), .A2(n_0_777), .B1(n_0_783), .B2(n_0_745), 
      .C1(n_0_781), .C2(n_0_714), .ZN(n_0_33_28));
   INV_X1 i_0_33_57 (.A(n_0_33_28), .ZN(n_0_811));
   AOI222_X1 i_0_33_58 (.A1(n_0_782), .A2(n_0_778), .B1(n_0_783), .B2(n_0_746), 
      .C1(n_0_781), .C2(n_0_715), .ZN(n_0_33_29));
   INV_X1 i_0_33_59 (.A(n_0_33_29), .ZN(n_0_812));
   AND2_X1 i_0_33_60 (.A1(n_0_781), .A2(n_0_716), .ZN(n_0_33_30));
   AOI221_X1 i_0_33_61 (.A(n_0_33_30), .B1(n_0_782), .B2(n_0_779), .C1(n_0_783), 
      .C2(n_0_747), .ZN(n_0_33_31));
   INV_X1 i_0_33_62 (.A(n_0_33_31), .ZN(n_0_813));
   AOI221_X1 i_0_33_63 (.A(n_0_33_30), .B1(n_0_782), .B2(n_0_780), .C1(n_0_783), 
      .C2(n_0_748), .ZN(n_0_33_32));
   INV_X1 i_0_33_64 (.A(n_0_33_32), .ZN(n_0_814));
   datapath__0_32 i_0_34 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_17, 
      n_0_814, n_0_813, n_0_812, n_0_811, n_0_810, n_0_809, n_0_808, n_0_807, 
      n_0_806, n_0_805, n_0_804, n_0_803, n_0_802, n_0_801, n_0_800, n_0_799, 
      n_0_798, n_0_797, n_0_796, n_0_795, n_0_794, n_0_793, n_0_792, n_0_791, 
      n_0_790, n_0_789, n_0_788, n_0_787, n_0_786, n_0_785, n_0_784}), .p_2({
      n_0_846, n_0_845, n_0_844, n_0_843, n_0_842, n_0_841, n_0_840, n_0_839, 
      n_0_838, n_0_837, n_0_836, n_0_835, n_0_834, n_0_833, n_0_832, n_0_831, 
      n_0_830, n_0_829, n_0_828, n_0_827, n_0_826, n_0_825, n_0_824, n_0_823, 
      n_0_822, n_0_821, n_0_820, n_0_819, n_0_818, n_0_817, n_0_816, n_0_815}));
   datapath__0_33 i_0_35 (.multiplicand2(multiplicand2), .p_0({uc_18, n_0_814, 
      n_0_813, n_0_812, n_0_811, n_0_810, n_0_809, n_0_808, n_0_807, n_0_806, 
      n_0_805, n_0_804, n_0_803, n_0_802, n_0_801, n_0_800, n_0_799, n_0_798, 
      n_0_797, n_0_796, n_0_795, n_0_794, n_0_793, n_0_792, n_0_791, n_0_790, 
      n_0_789, n_0_788, n_0_787, n_0_786, n_0_785, n_0_784}), .p_1({n_0_878, 
      n_0_877, n_0_876, n_0_875, n_0_874, n_0_873, n_0_872, n_0_871, n_0_870, 
      n_0_869, n_0_868, n_0_867, n_0_866, n_0_865, n_0_864, n_0_863, n_0_862, 
      n_0_861, n_0_860, n_0_859, n_0_858, n_0_857, n_0_856, n_0_855, n_0_854, 
      n_0_853, n_0_852, n_0_851, n_0_850, n_0_849, n_0_848, n_0_847}));
   INV_X1 i_0_36_0 (.A(multiplier2[9]), .ZN(n_0_36_0));
   AND2_X1 i_0_36_1 (.A1(n_0_36_0), .A2(multiplier2[8]), .ZN(n_0_880));
   NOR2_X1 i_0_36_2 (.A1(n_0_36_0), .A2(multiplier2[8]), .ZN(n_0_881));
   NOR2_X1 i_0_36_3 (.A1(n_0_880), .A2(n_0_881), .ZN(n_0_879));
   AOI222_X1 i_0_37_0 (.A1(n_0_847), .A2(n_0_880), .B1(n_0_815), .B2(n_0_881), 
      .C1(n_0_784), .C2(n_0_879), .ZN(n_0_37_0));
   INV_X1 i_0_37_1 (.A(n_0_37_0), .ZN(product[9]));
   AOI222_X1 i_0_37_2 (.A1(n_0_880), .A2(n_0_848), .B1(n_0_881), .B2(n_0_816), 
      .C1(n_0_879), .C2(n_0_785), .ZN(n_0_37_1));
   INV_X1 i_0_37_3 (.A(n_0_37_1), .ZN(n_0_882));
   AOI222_X1 i_0_37_4 (.A1(n_0_880), .A2(n_0_849), .B1(n_0_881), .B2(n_0_817), 
      .C1(n_0_879), .C2(n_0_786), .ZN(n_0_37_2));
   INV_X1 i_0_37_5 (.A(n_0_37_2), .ZN(n_0_883));
   AOI222_X1 i_0_37_6 (.A1(n_0_880), .A2(n_0_850), .B1(n_0_881), .B2(n_0_818), 
      .C1(n_0_879), .C2(n_0_787), .ZN(n_0_37_3));
   INV_X1 i_0_37_7 (.A(n_0_37_3), .ZN(n_0_884));
   AOI222_X1 i_0_37_8 (.A1(n_0_880), .A2(n_0_851), .B1(n_0_881), .B2(n_0_819), 
      .C1(n_0_879), .C2(n_0_788), .ZN(n_0_37_4));
   INV_X1 i_0_37_9 (.A(n_0_37_4), .ZN(n_0_885));
   AOI222_X1 i_0_37_10 (.A1(n_0_880), .A2(n_0_852), .B1(n_0_881), .B2(n_0_820), 
      .C1(n_0_879), .C2(n_0_789), .ZN(n_0_37_5));
   INV_X1 i_0_37_11 (.A(n_0_37_5), .ZN(n_0_886));
   AOI222_X1 i_0_37_12 (.A1(n_0_880), .A2(n_0_853), .B1(n_0_881), .B2(n_0_821), 
      .C1(n_0_879), .C2(n_0_790), .ZN(n_0_37_6));
   INV_X1 i_0_37_13 (.A(n_0_37_6), .ZN(n_0_887));
   AOI222_X1 i_0_37_14 (.A1(n_0_880), .A2(n_0_854), .B1(n_0_881), .B2(n_0_822), 
      .C1(n_0_879), .C2(n_0_791), .ZN(n_0_37_7));
   INV_X1 i_0_37_15 (.A(n_0_37_7), .ZN(n_0_888));
   AOI222_X1 i_0_37_16 (.A1(n_0_880), .A2(n_0_855), .B1(n_0_881), .B2(n_0_823), 
      .C1(n_0_879), .C2(n_0_792), .ZN(n_0_37_8));
   INV_X1 i_0_37_17 (.A(n_0_37_8), .ZN(n_0_889));
   AOI222_X1 i_0_37_18 (.A1(n_0_880), .A2(n_0_856), .B1(n_0_881), .B2(n_0_824), 
      .C1(n_0_879), .C2(n_0_793), .ZN(n_0_37_9));
   INV_X1 i_0_37_19 (.A(n_0_37_9), .ZN(n_0_890));
   AOI222_X1 i_0_37_20 (.A1(n_0_880), .A2(n_0_857), .B1(n_0_881), .B2(n_0_825), 
      .C1(n_0_879), .C2(n_0_794), .ZN(n_0_37_10));
   INV_X1 i_0_37_21 (.A(n_0_37_10), .ZN(n_0_891));
   AOI222_X1 i_0_37_22 (.A1(n_0_880), .A2(n_0_858), .B1(n_0_881), .B2(n_0_826), 
      .C1(n_0_879), .C2(n_0_795), .ZN(n_0_37_11));
   INV_X1 i_0_37_23 (.A(n_0_37_11), .ZN(n_0_892));
   AOI222_X1 i_0_37_24 (.A1(n_0_880), .A2(n_0_859), .B1(n_0_881), .B2(n_0_827), 
      .C1(n_0_879), .C2(n_0_796), .ZN(n_0_37_12));
   INV_X1 i_0_37_25 (.A(n_0_37_12), .ZN(n_0_893));
   AOI222_X1 i_0_37_26 (.A1(n_0_880), .A2(n_0_860), .B1(n_0_881), .B2(n_0_828), 
      .C1(n_0_879), .C2(n_0_797), .ZN(n_0_37_13));
   INV_X1 i_0_37_27 (.A(n_0_37_13), .ZN(n_0_894));
   AOI222_X1 i_0_37_28 (.A1(n_0_880), .A2(n_0_861), .B1(n_0_881), .B2(n_0_829), 
      .C1(n_0_879), .C2(n_0_798), .ZN(n_0_37_14));
   INV_X1 i_0_37_29 (.A(n_0_37_14), .ZN(n_0_895));
   AOI222_X1 i_0_37_30 (.A1(n_0_880), .A2(n_0_862), .B1(n_0_881), .B2(n_0_830), 
      .C1(n_0_879), .C2(n_0_799), .ZN(n_0_37_15));
   INV_X1 i_0_37_31 (.A(n_0_37_15), .ZN(n_0_896));
   AOI222_X1 i_0_37_32 (.A1(n_0_880), .A2(n_0_863), .B1(n_0_881), .B2(n_0_831), 
      .C1(n_0_879), .C2(n_0_800), .ZN(n_0_37_16));
   INV_X1 i_0_37_33 (.A(n_0_37_16), .ZN(n_0_897));
   AOI222_X1 i_0_37_34 (.A1(n_0_880), .A2(n_0_864), .B1(n_0_881), .B2(n_0_832), 
      .C1(n_0_879), .C2(n_0_801), .ZN(n_0_37_17));
   INV_X1 i_0_37_35 (.A(n_0_37_17), .ZN(n_0_898));
   AOI222_X1 i_0_37_36 (.A1(n_0_880), .A2(n_0_865), .B1(n_0_881), .B2(n_0_833), 
      .C1(n_0_879), .C2(n_0_802), .ZN(n_0_37_18));
   INV_X1 i_0_37_37 (.A(n_0_37_18), .ZN(n_0_899));
   AOI222_X1 i_0_37_38 (.A1(n_0_880), .A2(n_0_866), .B1(n_0_881), .B2(n_0_834), 
      .C1(n_0_879), .C2(n_0_803), .ZN(n_0_37_19));
   INV_X1 i_0_37_39 (.A(n_0_37_19), .ZN(n_0_900));
   AOI222_X1 i_0_37_40 (.A1(n_0_880), .A2(n_0_867), .B1(n_0_881), .B2(n_0_835), 
      .C1(n_0_879), .C2(n_0_804), .ZN(n_0_37_20));
   INV_X1 i_0_37_41 (.A(n_0_37_20), .ZN(n_0_901));
   AOI222_X1 i_0_37_42 (.A1(n_0_880), .A2(n_0_868), .B1(n_0_881), .B2(n_0_836), 
      .C1(n_0_879), .C2(n_0_805), .ZN(n_0_37_21));
   INV_X1 i_0_37_43 (.A(n_0_37_21), .ZN(n_0_902));
   AOI222_X1 i_0_37_44 (.A1(n_0_880), .A2(n_0_869), .B1(n_0_881), .B2(n_0_837), 
      .C1(n_0_879), .C2(n_0_806), .ZN(n_0_37_22));
   INV_X1 i_0_37_45 (.A(n_0_37_22), .ZN(n_0_903));
   AOI222_X1 i_0_37_46 (.A1(n_0_880), .A2(n_0_870), .B1(n_0_881), .B2(n_0_838), 
      .C1(n_0_879), .C2(n_0_807), .ZN(n_0_37_23));
   INV_X1 i_0_37_47 (.A(n_0_37_23), .ZN(n_0_904));
   AOI222_X1 i_0_37_48 (.A1(n_0_880), .A2(n_0_871), .B1(n_0_881), .B2(n_0_839), 
      .C1(n_0_879), .C2(n_0_808), .ZN(n_0_37_24));
   INV_X1 i_0_37_49 (.A(n_0_37_24), .ZN(n_0_905));
   AOI222_X1 i_0_37_50 (.A1(n_0_880), .A2(n_0_872), .B1(n_0_881), .B2(n_0_840), 
      .C1(n_0_879), .C2(n_0_809), .ZN(n_0_37_25));
   INV_X1 i_0_37_51 (.A(n_0_37_25), .ZN(n_0_906));
   AOI222_X1 i_0_37_52 (.A1(n_0_880), .A2(n_0_873), .B1(n_0_881), .B2(n_0_841), 
      .C1(n_0_879), .C2(n_0_810), .ZN(n_0_37_26));
   INV_X1 i_0_37_53 (.A(n_0_37_26), .ZN(n_0_907));
   AOI222_X1 i_0_37_54 (.A1(n_0_880), .A2(n_0_874), .B1(n_0_881), .B2(n_0_842), 
      .C1(n_0_879), .C2(n_0_811), .ZN(n_0_37_27));
   INV_X1 i_0_37_55 (.A(n_0_37_27), .ZN(n_0_908));
   AOI222_X1 i_0_37_56 (.A1(n_0_880), .A2(n_0_875), .B1(n_0_881), .B2(n_0_843), 
      .C1(n_0_879), .C2(n_0_812), .ZN(n_0_37_28));
   INV_X1 i_0_37_57 (.A(n_0_37_28), .ZN(n_0_909));
   AOI222_X1 i_0_37_58 (.A1(n_0_880), .A2(n_0_876), .B1(n_0_881), .B2(n_0_844), 
      .C1(n_0_879), .C2(n_0_813), .ZN(n_0_37_29));
   INV_X1 i_0_37_59 (.A(n_0_37_29), .ZN(n_0_910));
   AND2_X1 i_0_37_60 (.A1(n_0_879), .A2(n_0_814), .ZN(n_0_37_30));
   AOI221_X1 i_0_37_61 (.A(n_0_37_30), .B1(n_0_880), .B2(n_0_877), .C1(n_0_881), 
      .C2(n_0_845), .ZN(n_0_37_31));
   INV_X1 i_0_37_62 (.A(n_0_37_31), .ZN(n_0_911));
   AOI221_X1 i_0_37_63 (.A(n_0_37_30), .B1(n_0_880), .B2(n_0_878), .C1(n_0_881), 
      .C2(n_0_846), .ZN(n_0_37_32));
   INV_X1 i_0_37_64 (.A(n_0_37_32), .ZN(n_0_912));
   datapath__0_36 i_0_38 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_19, 
      n_0_912, n_0_911, n_0_910, n_0_909, n_0_908, n_0_907, n_0_906, n_0_905, 
      n_0_904, n_0_903, n_0_902, n_0_901, n_0_900, n_0_899, n_0_898, n_0_897, 
      n_0_896, n_0_895, n_0_894, n_0_893, n_0_892, n_0_891, n_0_890, n_0_889, 
      n_0_888, n_0_887, n_0_886, n_0_885, n_0_884, n_0_883, n_0_882}), .p_2({
      n_0_944, n_0_943, n_0_942, n_0_941, n_0_940, n_0_939, n_0_938, n_0_937, 
      n_0_936, n_0_935, n_0_934, n_0_933, n_0_932, n_0_931, n_0_930, n_0_929, 
      n_0_928, n_0_927, n_0_926, n_0_925, n_0_924, n_0_923, n_0_922, n_0_921, 
      n_0_920, n_0_919, n_0_918, n_0_917, n_0_916, n_0_915, n_0_914, n_0_913}));
   datapath__0_37 i_0_39 (.multiplicand2(multiplicand2), .p_0({uc_20, n_0_912, 
      n_0_911, n_0_910, n_0_909, n_0_908, n_0_907, n_0_906, n_0_905, n_0_904, 
      n_0_903, n_0_902, n_0_901, n_0_900, n_0_899, n_0_898, n_0_897, n_0_896, 
      n_0_895, n_0_894, n_0_893, n_0_892, n_0_891, n_0_890, n_0_889, n_0_888, 
      n_0_887, n_0_886, n_0_885, n_0_884, n_0_883, n_0_882}), .p_1({n_0_976, 
      n_0_975, n_0_974, n_0_973, n_0_972, n_0_971, n_0_970, n_0_969, n_0_968, 
      n_0_967, n_0_966, n_0_965, n_0_964, n_0_963, n_0_962, n_0_961, n_0_960, 
      n_0_959, n_0_958, n_0_957, n_0_956, n_0_955, n_0_954, n_0_953, n_0_952, 
      n_0_951, n_0_950, n_0_949, n_0_948, n_0_947, n_0_946, n_0_945}));
   INV_X1 i_0_40_0 (.A(multiplier2[10]), .ZN(n_0_40_0));
   AND2_X1 i_0_40_1 (.A1(n_0_40_0), .A2(multiplier2[9]), .ZN(n_0_978));
   NOR2_X1 i_0_40_2 (.A1(n_0_40_0), .A2(multiplier2[9]), .ZN(n_0_979));
   NOR2_X1 i_0_40_3 (.A1(n_0_978), .A2(n_0_979), .ZN(n_0_977));
   AOI222_X1 i_0_41_0 (.A1(n_0_945), .A2(n_0_978), .B1(n_0_913), .B2(n_0_979), 
      .C1(n_0_882), .C2(n_0_977), .ZN(n_0_41_0));
   INV_X1 i_0_41_1 (.A(n_0_41_0), .ZN(product[10]));
   AOI222_X1 i_0_41_2 (.A1(n_0_978), .A2(n_0_946), .B1(n_0_979), .B2(n_0_914), 
      .C1(n_0_977), .C2(n_0_883), .ZN(n_0_41_1));
   INV_X1 i_0_41_3 (.A(n_0_41_1), .ZN(n_0_980));
   AOI222_X1 i_0_41_4 (.A1(n_0_978), .A2(n_0_947), .B1(n_0_979), .B2(n_0_915), 
      .C1(n_0_977), .C2(n_0_884), .ZN(n_0_41_2));
   INV_X1 i_0_41_5 (.A(n_0_41_2), .ZN(n_0_981));
   AOI222_X1 i_0_41_6 (.A1(n_0_978), .A2(n_0_948), .B1(n_0_979), .B2(n_0_916), 
      .C1(n_0_977), .C2(n_0_885), .ZN(n_0_41_3));
   INV_X1 i_0_41_7 (.A(n_0_41_3), .ZN(n_0_982));
   AOI222_X1 i_0_41_8 (.A1(n_0_978), .A2(n_0_949), .B1(n_0_979), .B2(n_0_917), 
      .C1(n_0_977), .C2(n_0_886), .ZN(n_0_41_4));
   INV_X1 i_0_41_9 (.A(n_0_41_4), .ZN(n_0_983));
   AOI222_X1 i_0_41_10 (.A1(n_0_978), .A2(n_0_950), .B1(n_0_979), .B2(n_0_918), 
      .C1(n_0_977), .C2(n_0_887), .ZN(n_0_41_5));
   INV_X1 i_0_41_11 (.A(n_0_41_5), .ZN(n_0_984));
   AOI222_X1 i_0_41_12 (.A1(n_0_978), .A2(n_0_951), .B1(n_0_979), .B2(n_0_919), 
      .C1(n_0_977), .C2(n_0_888), .ZN(n_0_41_6));
   INV_X1 i_0_41_13 (.A(n_0_41_6), .ZN(n_0_985));
   AOI222_X1 i_0_41_14 (.A1(n_0_978), .A2(n_0_952), .B1(n_0_979), .B2(n_0_920), 
      .C1(n_0_977), .C2(n_0_889), .ZN(n_0_41_7));
   INV_X1 i_0_41_15 (.A(n_0_41_7), .ZN(n_0_986));
   AOI222_X1 i_0_41_16 (.A1(n_0_978), .A2(n_0_953), .B1(n_0_979), .B2(n_0_921), 
      .C1(n_0_977), .C2(n_0_890), .ZN(n_0_41_8));
   INV_X1 i_0_41_17 (.A(n_0_41_8), .ZN(n_0_987));
   AOI222_X1 i_0_41_18 (.A1(n_0_978), .A2(n_0_954), .B1(n_0_979), .B2(n_0_922), 
      .C1(n_0_977), .C2(n_0_891), .ZN(n_0_41_9));
   INV_X1 i_0_41_19 (.A(n_0_41_9), .ZN(n_0_988));
   AOI222_X1 i_0_41_20 (.A1(n_0_978), .A2(n_0_955), .B1(n_0_979), .B2(n_0_923), 
      .C1(n_0_977), .C2(n_0_892), .ZN(n_0_41_10));
   INV_X1 i_0_41_21 (.A(n_0_41_10), .ZN(n_0_989));
   AOI222_X1 i_0_41_22 (.A1(n_0_978), .A2(n_0_956), .B1(n_0_979), .B2(n_0_924), 
      .C1(n_0_977), .C2(n_0_893), .ZN(n_0_41_11));
   INV_X1 i_0_41_23 (.A(n_0_41_11), .ZN(n_0_990));
   AOI222_X1 i_0_41_24 (.A1(n_0_978), .A2(n_0_957), .B1(n_0_979), .B2(n_0_925), 
      .C1(n_0_977), .C2(n_0_894), .ZN(n_0_41_12));
   INV_X1 i_0_41_25 (.A(n_0_41_12), .ZN(n_0_991));
   AOI222_X1 i_0_41_26 (.A1(n_0_978), .A2(n_0_958), .B1(n_0_979), .B2(n_0_926), 
      .C1(n_0_977), .C2(n_0_895), .ZN(n_0_41_13));
   INV_X1 i_0_41_27 (.A(n_0_41_13), .ZN(n_0_992));
   AOI222_X1 i_0_41_28 (.A1(n_0_978), .A2(n_0_959), .B1(n_0_979), .B2(n_0_927), 
      .C1(n_0_977), .C2(n_0_896), .ZN(n_0_41_14));
   INV_X1 i_0_41_29 (.A(n_0_41_14), .ZN(n_0_993));
   AOI222_X1 i_0_41_30 (.A1(n_0_978), .A2(n_0_960), .B1(n_0_979), .B2(n_0_928), 
      .C1(n_0_977), .C2(n_0_897), .ZN(n_0_41_15));
   INV_X1 i_0_41_31 (.A(n_0_41_15), .ZN(n_0_994));
   AOI222_X1 i_0_41_32 (.A1(n_0_978), .A2(n_0_961), .B1(n_0_979), .B2(n_0_929), 
      .C1(n_0_977), .C2(n_0_898), .ZN(n_0_41_16));
   INV_X1 i_0_41_33 (.A(n_0_41_16), .ZN(n_0_995));
   AOI222_X1 i_0_41_34 (.A1(n_0_978), .A2(n_0_962), .B1(n_0_979), .B2(n_0_930), 
      .C1(n_0_977), .C2(n_0_899), .ZN(n_0_41_17));
   INV_X1 i_0_41_35 (.A(n_0_41_17), .ZN(n_0_996));
   AOI222_X1 i_0_41_36 (.A1(n_0_978), .A2(n_0_963), .B1(n_0_979), .B2(n_0_931), 
      .C1(n_0_977), .C2(n_0_900), .ZN(n_0_41_18));
   INV_X1 i_0_41_37 (.A(n_0_41_18), .ZN(n_0_997));
   AOI222_X1 i_0_41_38 (.A1(n_0_978), .A2(n_0_964), .B1(n_0_979), .B2(n_0_932), 
      .C1(n_0_977), .C2(n_0_901), .ZN(n_0_41_19));
   INV_X1 i_0_41_39 (.A(n_0_41_19), .ZN(n_0_998));
   AOI222_X1 i_0_41_40 (.A1(n_0_978), .A2(n_0_965), .B1(n_0_979), .B2(n_0_933), 
      .C1(n_0_977), .C2(n_0_902), .ZN(n_0_41_20));
   INV_X1 i_0_41_41 (.A(n_0_41_20), .ZN(n_0_999));
   AOI222_X1 i_0_41_42 (.A1(n_0_978), .A2(n_0_966), .B1(n_0_979), .B2(n_0_934), 
      .C1(n_0_977), .C2(n_0_903), .ZN(n_0_41_21));
   INV_X1 i_0_41_43 (.A(n_0_41_21), .ZN(n_0_1000));
   AOI222_X1 i_0_41_44 (.A1(n_0_978), .A2(n_0_967), .B1(n_0_979), .B2(n_0_935), 
      .C1(n_0_977), .C2(n_0_904), .ZN(n_0_41_22));
   INV_X1 i_0_41_45 (.A(n_0_41_22), .ZN(n_0_1001));
   AOI222_X1 i_0_41_46 (.A1(n_0_978), .A2(n_0_968), .B1(n_0_979), .B2(n_0_936), 
      .C1(n_0_977), .C2(n_0_905), .ZN(n_0_41_23));
   INV_X1 i_0_41_47 (.A(n_0_41_23), .ZN(n_0_1002));
   AOI222_X1 i_0_41_48 (.A1(n_0_978), .A2(n_0_969), .B1(n_0_979), .B2(n_0_937), 
      .C1(n_0_977), .C2(n_0_906), .ZN(n_0_41_24));
   INV_X1 i_0_41_49 (.A(n_0_41_24), .ZN(n_0_1003));
   AOI222_X1 i_0_41_50 (.A1(n_0_978), .A2(n_0_970), .B1(n_0_979), .B2(n_0_938), 
      .C1(n_0_977), .C2(n_0_907), .ZN(n_0_41_25));
   INV_X1 i_0_41_51 (.A(n_0_41_25), .ZN(n_0_1004));
   AOI222_X1 i_0_41_52 (.A1(n_0_978), .A2(n_0_971), .B1(n_0_979), .B2(n_0_939), 
      .C1(n_0_977), .C2(n_0_908), .ZN(n_0_41_26));
   INV_X1 i_0_41_53 (.A(n_0_41_26), .ZN(n_0_1005));
   AOI222_X1 i_0_41_54 (.A1(n_0_978), .A2(n_0_972), .B1(n_0_979), .B2(n_0_940), 
      .C1(n_0_977), .C2(n_0_909), .ZN(n_0_41_27));
   INV_X1 i_0_41_55 (.A(n_0_41_27), .ZN(n_0_1006));
   AOI222_X1 i_0_41_56 (.A1(n_0_978), .A2(n_0_973), .B1(n_0_979), .B2(n_0_941), 
      .C1(n_0_977), .C2(n_0_910), .ZN(n_0_41_28));
   INV_X1 i_0_41_57 (.A(n_0_41_28), .ZN(n_0_1007));
   AOI222_X1 i_0_41_58 (.A1(n_0_978), .A2(n_0_974), .B1(n_0_979), .B2(n_0_942), 
      .C1(n_0_977), .C2(n_0_911), .ZN(n_0_41_29));
   INV_X1 i_0_41_59 (.A(n_0_41_29), .ZN(n_0_1008));
   AND2_X1 i_0_41_60 (.A1(n_0_977), .A2(n_0_912), .ZN(n_0_41_30));
   AOI221_X1 i_0_41_61 (.A(n_0_41_30), .B1(n_0_978), .B2(n_0_975), .C1(n_0_979), 
      .C2(n_0_943), .ZN(n_0_41_31));
   INV_X1 i_0_41_62 (.A(n_0_41_31), .ZN(n_0_1009));
   AOI221_X1 i_0_41_63 (.A(n_0_41_30), .B1(n_0_978), .B2(n_0_976), .C1(n_0_979), 
      .C2(n_0_944), .ZN(n_0_41_32));
   INV_X1 i_0_41_64 (.A(n_0_41_32), .ZN(n_0_1010));
   datapath__0_40 i_0_42 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_21, 
      n_0_1010, n_0_1009, n_0_1008, n_0_1007, n_0_1006, n_0_1005, n_0_1004, 
      n_0_1003, n_0_1002, n_0_1001, n_0_1000, n_0_999, n_0_998, n_0_997, n_0_996, 
      n_0_995, n_0_994, n_0_993, n_0_992, n_0_991, n_0_990, n_0_989, n_0_988, 
      n_0_987, n_0_986, n_0_985, n_0_984, n_0_983, n_0_982, n_0_981, n_0_980}), 
      .p_2({n_0_1042, n_0_1041, n_0_1040, n_0_1039, n_0_1038, n_0_1037, n_0_1036, 
      n_0_1035, n_0_1034, n_0_1033, n_0_1032, n_0_1031, n_0_1030, n_0_1029, 
      n_0_1028, n_0_1027, n_0_1026, n_0_1025, n_0_1024, n_0_1023, n_0_1022, 
      n_0_1021, n_0_1020, n_0_1019, n_0_1018, n_0_1017, n_0_1016, n_0_1015, 
      n_0_1014, n_0_1013, n_0_1012, n_0_1011}));
   datapath__0_41 i_0_43 (.multiplicand2(multiplicand2), .p_0({uc_22, n_0_1010, 
      n_0_1009, n_0_1008, n_0_1007, n_0_1006, n_0_1005, n_0_1004, n_0_1003, 
      n_0_1002, n_0_1001, n_0_1000, n_0_999, n_0_998, n_0_997, n_0_996, n_0_995, 
      n_0_994, n_0_993, n_0_992, n_0_991, n_0_990, n_0_989, n_0_988, n_0_987, 
      n_0_986, n_0_985, n_0_984, n_0_983, n_0_982, n_0_981, n_0_980}), .p_1({
      n_0_1074, n_0_1073, n_0_1072, n_0_1071, n_0_1070, n_0_1069, n_0_1068, 
      n_0_1067, n_0_1066, n_0_1065, n_0_1064, n_0_1063, n_0_1062, n_0_1061, 
      n_0_1060, n_0_1059, n_0_1058, n_0_1057, n_0_1056, n_0_1055, n_0_1054, 
      n_0_1053, n_0_1052, n_0_1051, n_0_1050, n_0_1049, n_0_1048, n_0_1047, 
      n_0_1046, n_0_1045, n_0_1044, n_0_1043}));
   INV_X1 i_0_44_0 (.A(multiplier2[11]), .ZN(n_0_44_0));
   AND2_X1 i_0_44_1 (.A1(n_0_44_0), .A2(multiplier2[10]), .ZN(n_0_1076));
   NOR2_X1 i_0_44_2 (.A1(n_0_44_0), .A2(multiplier2[10]), .ZN(n_0_1077));
   NOR2_X1 i_0_44_3 (.A1(n_0_1076), .A2(n_0_1077), .ZN(n_0_1075));
   AOI222_X1 i_0_45_0 (.A1(n_0_1043), .A2(n_0_1076), .B1(n_0_1011), .B2(n_0_1077), 
      .C1(n_0_980), .C2(n_0_1075), .ZN(n_0_45_0));
   INV_X1 i_0_45_1 (.A(n_0_45_0), .ZN(product[11]));
   AOI222_X1 i_0_45_2 (.A1(n_0_1076), .A2(n_0_1044), .B1(n_0_1077), .B2(n_0_1012), 
      .C1(n_0_1075), .C2(n_0_981), .ZN(n_0_45_1));
   INV_X1 i_0_45_3 (.A(n_0_45_1), .ZN(n_0_1078));
   AOI222_X1 i_0_45_4 (.A1(n_0_1076), .A2(n_0_1045), .B1(n_0_1077), .B2(n_0_1013), 
      .C1(n_0_1075), .C2(n_0_982), .ZN(n_0_45_2));
   INV_X1 i_0_45_5 (.A(n_0_45_2), .ZN(n_0_1079));
   AOI222_X1 i_0_45_6 (.A1(n_0_1076), .A2(n_0_1046), .B1(n_0_1077), .B2(n_0_1014), 
      .C1(n_0_1075), .C2(n_0_983), .ZN(n_0_45_3));
   INV_X1 i_0_45_7 (.A(n_0_45_3), .ZN(n_0_1080));
   AOI222_X1 i_0_45_8 (.A1(n_0_1076), .A2(n_0_1047), .B1(n_0_1077), .B2(n_0_1015), 
      .C1(n_0_1075), .C2(n_0_984), .ZN(n_0_45_4));
   INV_X1 i_0_45_9 (.A(n_0_45_4), .ZN(n_0_1081));
   AOI222_X1 i_0_45_10 (.A1(n_0_1076), .A2(n_0_1048), .B1(n_0_1077), .B2(
      n_0_1016), .C1(n_0_1075), .C2(n_0_985), .ZN(n_0_45_5));
   INV_X1 i_0_45_11 (.A(n_0_45_5), .ZN(n_0_1082));
   AOI222_X1 i_0_45_12 (.A1(n_0_1076), .A2(n_0_1049), .B1(n_0_1077), .B2(
      n_0_1017), .C1(n_0_1075), .C2(n_0_986), .ZN(n_0_45_6));
   INV_X1 i_0_45_13 (.A(n_0_45_6), .ZN(n_0_1083));
   AOI222_X1 i_0_45_14 (.A1(n_0_1076), .A2(n_0_1050), .B1(n_0_1077), .B2(
      n_0_1018), .C1(n_0_1075), .C2(n_0_987), .ZN(n_0_45_7));
   INV_X1 i_0_45_15 (.A(n_0_45_7), .ZN(n_0_1084));
   AOI222_X1 i_0_45_16 (.A1(n_0_1076), .A2(n_0_1051), .B1(n_0_1077), .B2(
      n_0_1019), .C1(n_0_1075), .C2(n_0_988), .ZN(n_0_45_8));
   INV_X1 i_0_45_17 (.A(n_0_45_8), .ZN(n_0_1085));
   AOI222_X1 i_0_45_18 (.A1(n_0_1076), .A2(n_0_1052), .B1(n_0_1077), .B2(
      n_0_1020), .C1(n_0_1075), .C2(n_0_989), .ZN(n_0_45_9));
   INV_X1 i_0_45_19 (.A(n_0_45_9), .ZN(n_0_1086));
   AOI222_X1 i_0_45_20 (.A1(n_0_1076), .A2(n_0_1053), .B1(n_0_1077), .B2(
      n_0_1021), .C1(n_0_1075), .C2(n_0_990), .ZN(n_0_45_10));
   INV_X1 i_0_45_21 (.A(n_0_45_10), .ZN(n_0_1087));
   AOI222_X1 i_0_45_22 (.A1(n_0_1076), .A2(n_0_1054), .B1(n_0_1077), .B2(
      n_0_1022), .C1(n_0_1075), .C2(n_0_991), .ZN(n_0_45_11));
   INV_X1 i_0_45_23 (.A(n_0_45_11), .ZN(n_0_1088));
   AOI222_X1 i_0_45_24 (.A1(n_0_1076), .A2(n_0_1055), .B1(n_0_1077), .B2(
      n_0_1023), .C1(n_0_1075), .C2(n_0_992), .ZN(n_0_45_12));
   INV_X1 i_0_45_25 (.A(n_0_45_12), .ZN(n_0_1089));
   AOI222_X1 i_0_45_26 (.A1(n_0_1076), .A2(n_0_1056), .B1(n_0_1077), .B2(
      n_0_1024), .C1(n_0_1075), .C2(n_0_993), .ZN(n_0_45_13));
   INV_X1 i_0_45_27 (.A(n_0_45_13), .ZN(n_0_1090));
   AOI222_X1 i_0_45_28 (.A1(n_0_1076), .A2(n_0_1057), .B1(n_0_1077), .B2(
      n_0_1025), .C1(n_0_1075), .C2(n_0_994), .ZN(n_0_45_14));
   INV_X1 i_0_45_29 (.A(n_0_45_14), .ZN(n_0_1091));
   AOI222_X1 i_0_45_30 (.A1(n_0_1076), .A2(n_0_1058), .B1(n_0_1077), .B2(
      n_0_1026), .C1(n_0_1075), .C2(n_0_995), .ZN(n_0_45_15));
   INV_X1 i_0_45_31 (.A(n_0_45_15), .ZN(n_0_1092));
   AOI222_X1 i_0_45_32 (.A1(n_0_1076), .A2(n_0_1059), .B1(n_0_1077), .B2(
      n_0_1027), .C1(n_0_1075), .C2(n_0_996), .ZN(n_0_45_16));
   INV_X1 i_0_45_33 (.A(n_0_45_16), .ZN(n_0_1093));
   AOI222_X1 i_0_45_34 (.A1(n_0_1076), .A2(n_0_1060), .B1(n_0_1077), .B2(
      n_0_1028), .C1(n_0_1075), .C2(n_0_997), .ZN(n_0_45_17));
   INV_X1 i_0_45_35 (.A(n_0_45_17), .ZN(n_0_1094));
   AOI222_X1 i_0_45_36 (.A1(n_0_1076), .A2(n_0_1061), .B1(n_0_1077), .B2(
      n_0_1029), .C1(n_0_1075), .C2(n_0_998), .ZN(n_0_45_18));
   INV_X1 i_0_45_37 (.A(n_0_45_18), .ZN(n_0_1095));
   AOI222_X1 i_0_45_38 (.A1(n_0_1076), .A2(n_0_1062), .B1(n_0_1077), .B2(
      n_0_1030), .C1(n_0_1075), .C2(n_0_999), .ZN(n_0_45_19));
   INV_X1 i_0_45_39 (.A(n_0_45_19), .ZN(n_0_1096));
   AOI222_X1 i_0_45_40 (.A1(n_0_1076), .A2(n_0_1063), .B1(n_0_1077), .B2(
      n_0_1031), .C1(n_0_1075), .C2(n_0_1000), .ZN(n_0_45_20));
   INV_X1 i_0_45_41 (.A(n_0_45_20), .ZN(n_0_1097));
   AOI222_X1 i_0_45_42 (.A1(n_0_1076), .A2(n_0_1064), .B1(n_0_1077), .B2(
      n_0_1032), .C1(n_0_1075), .C2(n_0_1001), .ZN(n_0_45_21));
   INV_X1 i_0_45_43 (.A(n_0_45_21), .ZN(n_0_1098));
   AOI222_X1 i_0_45_44 (.A1(n_0_1076), .A2(n_0_1065), .B1(n_0_1077), .B2(
      n_0_1033), .C1(n_0_1075), .C2(n_0_1002), .ZN(n_0_45_22));
   INV_X1 i_0_45_45 (.A(n_0_45_22), .ZN(n_0_1099));
   AOI222_X1 i_0_45_46 (.A1(n_0_1076), .A2(n_0_1066), .B1(n_0_1077), .B2(
      n_0_1034), .C1(n_0_1075), .C2(n_0_1003), .ZN(n_0_45_23));
   INV_X1 i_0_45_47 (.A(n_0_45_23), .ZN(n_0_1100));
   AOI222_X1 i_0_45_48 (.A1(n_0_1076), .A2(n_0_1067), .B1(n_0_1077), .B2(
      n_0_1035), .C1(n_0_1075), .C2(n_0_1004), .ZN(n_0_45_24));
   INV_X1 i_0_45_49 (.A(n_0_45_24), .ZN(n_0_1101));
   AOI222_X1 i_0_45_50 (.A1(n_0_1076), .A2(n_0_1068), .B1(n_0_1077), .B2(
      n_0_1036), .C1(n_0_1075), .C2(n_0_1005), .ZN(n_0_45_25));
   INV_X1 i_0_45_51 (.A(n_0_45_25), .ZN(n_0_1102));
   AOI222_X1 i_0_45_52 (.A1(n_0_1076), .A2(n_0_1069), .B1(n_0_1077), .B2(
      n_0_1037), .C1(n_0_1075), .C2(n_0_1006), .ZN(n_0_45_26));
   INV_X1 i_0_45_53 (.A(n_0_45_26), .ZN(n_0_1103));
   AOI222_X1 i_0_45_54 (.A1(n_0_1076), .A2(n_0_1070), .B1(n_0_1077), .B2(
      n_0_1038), .C1(n_0_1075), .C2(n_0_1007), .ZN(n_0_45_27));
   INV_X1 i_0_45_55 (.A(n_0_45_27), .ZN(n_0_1104));
   AOI222_X1 i_0_45_56 (.A1(n_0_1076), .A2(n_0_1071), .B1(n_0_1077), .B2(
      n_0_1039), .C1(n_0_1075), .C2(n_0_1008), .ZN(n_0_45_28));
   INV_X1 i_0_45_57 (.A(n_0_45_28), .ZN(n_0_1105));
   AOI222_X1 i_0_45_58 (.A1(n_0_1076), .A2(n_0_1072), .B1(n_0_1077), .B2(
      n_0_1040), .C1(n_0_1075), .C2(n_0_1009), .ZN(n_0_45_29));
   INV_X1 i_0_45_59 (.A(n_0_45_29), .ZN(n_0_1106));
   AND2_X1 i_0_45_60 (.A1(n_0_1075), .A2(n_0_1010), .ZN(n_0_45_30));
   AOI221_X1 i_0_45_61 (.A(n_0_45_30), .B1(n_0_1076), .B2(n_0_1073), .C1(
      n_0_1077), .C2(n_0_1041), .ZN(n_0_45_31));
   INV_X1 i_0_45_62 (.A(n_0_45_31), .ZN(n_0_1107));
   AOI221_X1 i_0_45_63 (.A(n_0_45_30), .B1(n_0_1076), .B2(n_0_1074), .C1(
      n_0_1077), .C2(n_0_1042), .ZN(n_0_45_32));
   INV_X1 i_0_45_64 (.A(n_0_45_32), .ZN(n_0_1108));
   datapath__0_44 i_0_46 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_23, 
      n_0_1108, n_0_1107, n_0_1106, n_0_1105, n_0_1104, n_0_1103, n_0_1102, 
      n_0_1101, n_0_1100, n_0_1099, n_0_1098, n_0_1097, n_0_1096, n_0_1095, 
      n_0_1094, n_0_1093, n_0_1092, n_0_1091, n_0_1090, n_0_1089, n_0_1088, 
      n_0_1087, n_0_1086, n_0_1085, n_0_1084, n_0_1083, n_0_1082, n_0_1081, 
      n_0_1080, n_0_1079, n_0_1078}), .p_2({n_0_1140, n_0_1139, n_0_1138, 
      n_0_1137, n_0_1136, n_0_1135, n_0_1134, n_0_1133, n_0_1132, n_0_1131, 
      n_0_1130, n_0_1129, n_0_1128, n_0_1127, n_0_1126, n_0_1125, n_0_1124, 
      n_0_1123, n_0_1122, n_0_1121, n_0_1120, n_0_1119, n_0_1118, n_0_1117, 
      n_0_1116, n_0_1115, n_0_1114, n_0_1113, n_0_1112, n_0_1111, n_0_1110, 
      n_0_1109}));
   datapath__0_45 i_0_47 (.multiplicand2(multiplicand2), .p_0({uc_24, n_0_1108, 
      n_0_1107, n_0_1106, n_0_1105, n_0_1104, n_0_1103, n_0_1102, n_0_1101, 
      n_0_1100, n_0_1099, n_0_1098, n_0_1097, n_0_1096, n_0_1095, n_0_1094, 
      n_0_1093, n_0_1092, n_0_1091, n_0_1090, n_0_1089, n_0_1088, n_0_1087, 
      n_0_1086, n_0_1085, n_0_1084, n_0_1083, n_0_1082, n_0_1081, n_0_1080, 
      n_0_1079, n_0_1078}), .p_1({n_0_1172, n_0_1171, n_0_1170, n_0_1169, 
      n_0_1168, n_0_1167, n_0_1166, n_0_1165, n_0_1164, n_0_1163, n_0_1162, 
      n_0_1161, n_0_1160, n_0_1159, n_0_1158, n_0_1157, n_0_1156, n_0_1155, 
      n_0_1154, n_0_1153, n_0_1152, n_0_1151, n_0_1150, n_0_1149, n_0_1148, 
      n_0_1147, n_0_1146, n_0_1145, n_0_1144, n_0_1143, n_0_1142, n_0_1141}));
   INV_X1 i_0_48_0 (.A(multiplier2[12]), .ZN(n_0_48_0));
   AND2_X1 i_0_48_1 (.A1(n_0_48_0), .A2(multiplier2[11]), .ZN(n_0_1174));
   NOR2_X1 i_0_48_2 (.A1(n_0_48_0), .A2(multiplier2[11]), .ZN(n_0_1175));
   NOR2_X1 i_0_48_3 (.A1(n_0_1174), .A2(n_0_1175), .ZN(n_0_1173));
   AOI222_X1 i_0_49_0 (.A1(n_0_1141), .A2(n_0_1174), .B1(n_0_1109), .B2(n_0_1175), 
      .C1(n_0_1078), .C2(n_0_1173), .ZN(n_0_49_0));
   INV_X1 i_0_49_1 (.A(n_0_49_0), .ZN(product[12]));
   AOI222_X1 i_0_49_2 (.A1(n_0_1174), .A2(n_0_1142), .B1(n_0_1175), .B2(n_0_1110), 
      .C1(n_0_1173), .C2(n_0_1079), .ZN(n_0_49_1));
   INV_X1 i_0_49_3 (.A(n_0_49_1), .ZN(n_0_1176));
   AOI222_X1 i_0_49_4 (.A1(n_0_1174), .A2(n_0_1143), .B1(n_0_1175), .B2(n_0_1111), 
      .C1(n_0_1173), .C2(n_0_1080), .ZN(n_0_49_2));
   INV_X1 i_0_49_5 (.A(n_0_49_2), .ZN(n_0_1177));
   AOI222_X1 i_0_49_6 (.A1(n_0_1174), .A2(n_0_1144), .B1(n_0_1175), .B2(n_0_1112), 
      .C1(n_0_1173), .C2(n_0_1081), .ZN(n_0_49_3));
   INV_X1 i_0_49_7 (.A(n_0_49_3), .ZN(n_0_1178));
   AOI222_X1 i_0_49_8 (.A1(n_0_1174), .A2(n_0_1145), .B1(n_0_1175), .B2(n_0_1113), 
      .C1(n_0_1173), .C2(n_0_1082), .ZN(n_0_49_4));
   INV_X1 i_0_49_9 (.A(n_0_49_4), .ZN(n_0_1179));
   AOI222_X1 i_0_49_10 (.A1(n_0_1174), .A2(n_0_1146), .B1(n_0_1175), .B2(
      n_0_1114), .C1(n_0_1173), .C2(n_0_1083), .ZN(n_0_49_5));
   INV_X1 i_0_49_11 (.A(n_0_49_5), .ZN(n_0_1180));
   AOI222_X1 i_0_49_12 (.A1(n_0_1174), .A2(n_0_1147), .B1(n_0_1175), .B2(
      n_0_1115), .C1(n_0_1173), .C2(n_0_1084), .ZN(n_0_49_6));
   INV_X1 i_0_49_13 (.A(n_0_49_6), .ZN(n_0_1181));
   AOI222_X1 i_0_49_14 (.A1(n_0_1174), .A2(n_0_1148), .B1(n_0_1175), .B2(
      n_0_1116), .C1(n_0_1173), .C2(n_0_1085), .ZN(n_0_49_7));
   INV_X1 i_0_49_15 (.A(n_0_49_7), .ZN(n_0_1182));
   AOI222_X1 i_0_49_16 (.A1(n_0_1174), .A2(n_0_1149), .B1(n_0_1175), .B2(
      n_0_1117), .C1(n_0_1173), .C2(n_0_1086), .ZN(n_0_49_8));
   INV_X1 i_0_49_17 (.A(n_0_49_8), .ZN(n_0_1183));
   AOI222_X1 i_0_49_18 (.A1(n_0_1174), .A2(n_0_1150), .B1(n_0_1175), .B2(
      n_0_1118), .C1(n_0_1173), .C2(n_0_1087), .ZN(n_0_49_9));
   INV_X1 i_0_49_19 (.A(n_0_49_9), .ZN(n_0_1184));
   AOI222_X1 i_0_49_20 (.A1(n_0_1174), .A2(n_0_1151), .B1(n_0_1175), .B2(
      n_0_1119), .C1(n_0_1173), .C2(n_0_1088), .ZN(n_0_49_10));
   INV_X1 i_0_49_21 (.A(n_0_49_10), .ZN(n_0_1185));
   AOI222_X1 i_0_49_22 (.A1(n_0_1174), .A2(n_0_1152), .B1(n_0_1175), .B2(
      n_0_1120), .C1(n_0_1173), .C2(n_0_1089), .ZN(n_0_49_11));
   INV_X1 i_0_49_23 (.A(n_0_49_11), .ZN(n_0_1186));
   AOI222_X1 i_0_49_24 (.A1(n_0_1174), .A2(n_0_1153), .B1(n_0_1175), .B2(
      n_0_1121), .C1(n_0_1173), .C2(n_0_1090), .ZN(n_0_49_12));
   INV_X1 i_0_49_25 (.A(n_0_49_12), .ZN(n_0_1187));
   AOI222_X1 i_0_49_26 (.A1(n_0_1174), .A2(n_0_1154), .B1(n_0_1175), .B2(
      n_0_1122), .C1(n_0_1173), .C2(n_0_1091), .ZN(n_0_49_13));
   INV_X1 i_0_49_27 (.A(n_0_49_13), .ZN(n_0_1188));
   AOI222_X1 i_0_49_28 (.A1(n_0_1174), .A2(n_0_1155), .B1(n_0_1175), .B2(
      n_0_1123), .C1(n_0_1173), .C2(n_0_1092), .ZN(n_0_49_14));
   INV_X1 i_0_49_29 (.A(n_0_49_14), .ZN(n_0_1189));
   AOI222_X1 i_0_49_30 (.A1(n_0_1174), .A2(n_0_1156), .B1(n_0_1175), .B2(
      n_0_1124), .C1(n_0_1173), .C2(n_0_1093), .ZN(n_0_49_15));
   INV_X1 i_0_49_31 (.A(n_0_49_15), .ZN(n_0_1190));
   AOI222_X1 i_0_49_32 (.A1(n_0_1174), .A2(n_0_1157), .B1(n_0_1175), .B2(
      n_0_1125), .C1(n_0_1173), .C2(n_0_1094), .ZN(n_0_49_16));
   INV_X1 i_0_49_33 (.A(n_0_49_16), .ZN(n_0_1191));
   AOI222_X1 i_0_49_34 (.A1(n_0_1174), .A2(n_0_1158), .B1(n_0_1175), .B2(
      n_0_1126), .C1(n_0_1173), .C2(n_0_1095), .ZN(n_0_49_17));
   INV_X1 i_0_49_35 (.A(n_0_49_17), .ZN(n_0_1192));
   AOI222_X1 i_0_49_36 (.A1(n_0_1174), .A2(n_0_1159), .B1(n_0_1175), .B2(
      n_0_1127), .C1(n_0_1173), .C2(n_0_1096), .ZN(n_0_49_18));
   INV_X1 i_0_49_37 (.A(n_0_49_18), .ZN(n_0_1193));
   AOI222_X1 i_0_49_38 (.A1(n_0_1174), .A2(n_0_1160), .B1(n_0_1175), .B2(
      n_0_1128), .C1(n_0_1173), .C2(n_0_1097), .ZN(n_0_49_19));
   INV_X1 i_0_49_39 (.A(n_0_49_19), .ZN(n_0_1194));
   AOI222_X1 i_0_49_40 (.A1(n_0_1174), .A2(n_0_1161), .B1(n_0_1175), .B2(
      n_0_1129), .C1(n_0_1173), .C2(n_0_1098), .ZN(n_0_49_20));
   INV_X1 i_0_49_41 (.A(n_0_49_20), .ZN(n_0_1195));
   AOI222_X1 i_0_49_42 (.A1(n_0_1174), .A2(n_0_1162), .B1(n_0_1175), .B2(
      n_0_1130), .C1(n_0_1173), .C2(n_0_1099), .ZN(n_0_49_21));
   INV_X1 i_0_49_43 (.A(n_0_49_21), .ZN(n_0_1196));
   AOI222_X1 i_0_49_44 (.A1(n_0_1174), .A2(n_0_1163), .B1(n_0_1175), .B2(
      n_0_1131), .C1(n_0_1173), .C2(n_0_1100), .ZN(n_0_49_22));
   INV_X1 i_0_49_45 (.A(n_0_49_22), .ZN(n_0_1197));
   AOI222_X1 i_0_49_46 (.A1(n_0_1174), .A2(n_0_1164), .B1(n_0_1175), .B2(
      n_0_1132), .C1(n_0_1173), .C2(n_0_1101), .ZN(n_0_49_23));
   INV_X1 i_0_49_47 (.A(n_0_49_23), .ZN(n_0_1198));
   AOI222_X1 i_0_49_48 (.A1(n_0_1174), .A2(n_0_1165), .B1(n_0_1175), .B2(
      n_0_1133), .C1(n_0_1173), .C2(n_0_1102), .ZN(n_0_49_24));
   INV_X1 i_0_49_49 (.A(n_0_49_24), .ZN(n_0_1199));
   AOI222_X1 i_0_49_50 (.A1(n_0_1174), .A2(n_0_1166), .B1(n_0_1175), .B2(
      n_0_1134), .C1(n_0_1173), .C2(n_0_1103), .ZN(n_0_49_25));
   INV_X1 i_0_49_51 (.A(n_0_49_25), .ZN(n_0_1200));
   AOI222_X1 i_0_49_52 (.A1(n_0_1174), .A2(n_0_1167), .B1(n_0_1175), .B2(
      n_0_1135), .C1(n_0_1173), .C2(n_0_1104), .ZN(n_0_49_26));
   INV_X1 i_0_49_53 (.A(n_0_49_26), .ZN(n_0_1201));
   AOI222_X1 i_0_49_54 (.A1(n_0_1174), .A2(n_0_1168), .B1(n_0_1175), .B2(
      n_0_1136), .C1(n_0_1173), .C2(n_0_1105), .ZN(n_0_49_27));
   INV_X1 i_0_49_55 (.A(n_0_49_27), .ZN(n_0_1202));
   AOI222_X1 i_0_49_56 (.A1(n_0_1174), .A2(n_0_1169), .B1(n_0_1175), .B2(
      n_0_1137), .C1(n_0_1173), .C2(n_0_1106), .ZN(n_0_49_28));
   INV_X1 i_0_49_57 (.A(n_0_49_28), .ZN(n_0_1203));
   AOI222_X1 i_0_49_58 (.A1(n_0_1174), .A2(n_0_1170), .B1(n_0_1175), .B2(
      n_0_1138), .C1(n_0_1173), .C2(n_0_1107), .ZN(n_0_49_29));
   INV_X1 i_0_49_59 (.A(n_0_49_29), .ZN(n_0_1204));
   AND2_X1 i_0_49_60 (.A1(n_0_1173), .A2(n_0_1108), .ZN(n_0_49_30));
   AOI221_X1 i_0_49_61 (.A(n_0_49_30), .B1(n_0_1174), .B2(n_0_1171), .C1(
      n_0_1175), .C2(n_0_1139), .ZN(n_0_49_31));
   INV_X1 i_0_49_62 (.A(n_0_49_31), .ZN(n_0_1205));
   AOI221_X1 i_0_49_63 (.A(n_0_49_30), .B1(n_0_1174), .B2(n_0_1172), .C1(
      n_0_1175), .C2(n_0_1140), .ZN(n_0_49_32));
   INV_X1 i_0_49_64 (.A(n_0_49_32), .ZN(n_0_1206));
   datapath__0_48 i_0_50 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_25, 
      n_0_1206, n_0_1205, n_0_1204, n_0_1203, n_0_1202, n_0_1201, n_0_1200, 
      n_0_1199, n_0_1198, n_0_1197, n_0_1196, n_0_1195, n_0_1194, n_0_1193, 
      n_0_1192, n_0_1191, n_0_1190, n_0_1189, n_0_1188, n_0_1187, n_0_1186, 
      n_0_1185, n_0_1184, n_0_1183, n_0_1182, n_0_1181, n_0_1180, n_0_1179, 
      n_0_1178, n_0_1177, n_0_1176}), .p_2({n_0_1238, n_0_1237, n_0_1236, 
      n_0_1235, n_0_1234, n_0_1233, n_0_1232, n_0_1231, n_0_1230, n_0_1229, 
      n_0_1228, n_0_1227, n_0_1226, n_0_1225, n_0_1224, n_0_1223, n_0_1222, 
      n_0_1221, n_0_1220, n_0_1219, n_0_1218, n_0_1217, n_0_1216, n_0_1215, 
      n_0_1214, n_0_1213, n_0_1212, n_0_1211, n_0_1210, n_0_1209, n_0_1208, 
      n_0_1207}));
   datapath__0_49 i_0_51 (.multiplicand2(multiplicand2), .p_0({uc_26, n_0_1206, 
      n_0_1205, n_0_1204, n_0_1203, n_0_1202, n_0_1201, n_0_1200, n_0_1199, 
      n_0_1198, n_0_1197, n_0_1196, n_0_1195, n_0_1194, n_0_1193, n_0_1192, 
      n_0_1191, n_0_1190, n_0_1189, n_0_1188, n_0_1187, n_0_1186, n_0_1185, 
      n_0_1184, n_0_1183, n_0_1182, n_0_1181, n_0_1180, n_0_1179, n_0_1178, 
      n_0_1177, n_0_1176}), .p_1({n_0_1270, n_0_1269, n_0_1268, n_0_1267, 
      n_0_1266, n_0_1265, n_0_1264, n_0_1263, n_0_1262, n_0_1261, n_0_1260, 
      n_0_1259, n_0_1258, n_0_1257, n_0_1256, n_0_1255, n_0_1254, n_0_1253, 
      n_0_1252, n_0_1251, n_0_1250, n_0_1249, n_0_1248, n_0_1247, n_0_1246, 
      n_0_1245, n_0_1244, n_0_1243, n_0_1242, n_0_1241, n_0_1240, n_0_1239}));
   INV_X1 i_0_52_0 (.A(multiplier2[13]), .ZN(n_0_52_0));
   AND2_X1 i_0_52_1 (.A1(n_0_52_0), .A2(multiplier2[12]), .ZN(n_0_1272));
   NOR2_X1 i_0_52_2 (.A1(n_0_52_0), .A2(multiplier2[12]), .ZN(n_0_1273));
   NOR2_X1 i_0_52_3 (.A1(n_0_1272), .A2(n_0_1273), .ZN(n_0_1271));
   AOI222_X1 i_0_53_0 (.A1(n_0_1239), .A2(n_0_1272), .B1(n_0_1207), .B2(n_0_1273), 
      .C1(n_0_1176), .C2(n_0_1271), .ZN(n_0_53_0));
   INV_X1 i_0_53_1 (.A(n_0_53_0), .ZN(product[13]));
   AOI222_X1 i_0_53_2 (.A1(n_0_1272), .A2(n_0_1240), .B1(n_0_1273), .B2(n_0_1208), 
      .C1(n_0_1271), .C2(n_0_1177), .ZN(n_0_53_1));
   INV_X1 i_0_53_3 (.A(n_0_53_1), .ZN(n_0_1274));
   AOI222_X1 i_0_53_4 (.A1(n_0_1272), .A2(n_0_1241), .B1(n_0_1273), .B2(n_0_1209), 
      .C1(n_0_1271), .C2(n_0_1178), .ZN(n_0_53_2));
   INV_X1 i_0_53_5 (.A(n_0_53_2), .ZN(n_0_1275));
   AOI222_X1 i_0_53_6 (.A1(n_0_1272), .A2(n_0_1242), .B1(n_0_1273), .B2(n_0_1210), 
      .C1(n_0_1271), .C2(n_0_1179), .ZN(n_0_53_3));
   INV_X1 i_0_53_7 (.A(n_0_53_3), .ZN(n_0_1276));
   AOI222_X1 i_0_53_8 (.A1(n_0_1272), .A2(n_0_1243), .B1(n_0_1273), .B2(n_0_1211), 
      .C1(n_0_1271), .C2(n_0_1180), .ZN(n_0_53_4));
   INV_X1 i_0_53_9 (.A(n_0_53_4), .ZN(n_0_1277));
   AOI222_X1 i_0_53_10 (.A1(n_0_1272), .A2(n_0_1244), .B1(n_0_1273), .B2(
      n_0_1212), .C1(n_0_1271), .C2(n_0_1181), .ZN(n_0_53_5));
   INV_X1 i_0_53_11 (.A(n_0_53_5), .ZN(n_0_1278));
   AOI222_X1 i_0_53_12 (.A1(n_0_1272), .A2(n_0_1245), .B1(n_0_1273), .B2(
      n_0_1213), .C1(n_0_1271), .C2(n_0_1182), .ZN(n_0_53_6));
   INV_X1 i_0_53_13 (.A(n_0_53_6), .ZN(n_0_1279));
   AOI222_X1 i_0_53_14 (.A1(n_0_1272), .A2(n_0_1246), .B1(n_0_1273), .B2(
      n_0_1214), .C1(n_0_1271), .C2(n_0_1183), .ZN(n_0_53_7));
   INV_X1 i_0_53_15 (.A(n_0_53_7), .ZN(n_0_1280));
   AOI222_X1 i_0_53_16 (.A1(n_0_1272), .A2(n_0_1247), .B1(n_0_1273), .B2(
      n_0_1215), .C1(n_0_1271), .C2(n_0_1184), .ZN(n_0_53_8));
   INV_X1 i_0_53_17 (.A(n_0_53_8), .ZN(n_0_1281));
   AOI222_X1 i_0_53_18 (.A1(n_0_1272), .A2(n_0_1248), .B1(n_0_1273), .B2(
      n_0_1216), .C1(n_0_1271), .C2(n_0_1185), .ZN(n_0_53_9));
   INV_X1 i_0_53_19 (.A(n_0_53_9), .ZN(n_0_1282));
   AOI222_X1 i_0_53_20 (.A1(n_0_1272), .A2(n_0_1249), .B1(n_0_1273), .B2(
      n_0_1217), .C1(n_0_1271), .C2(n_0_1186), .ZN(n_0_53_10));
   INV_X1 i_0_53_21 (.A(n_0_53_10), .ZN(n_0_1283));
   AOI222_X1 i_0_53_22 (.A1(n_0_1272), .A2(n_0_1250), .B1(n_0_1273), .B2(
      n_0_1218), .C1(n_0_1271), .C2(n_0_1187), .ZN(n_0_53_11));
   INV_X1 i_0_53_23 (.A(n_0_53_11), .ZN(n_0_1284));
   AOI222_X1 i_0_53_24 (.A1(n_0_1272), .A2(n_0_1251), .B1(n_0_1273), .B2(
      n_0_1219), .C1(n_0_1271), .C2(n_0_1188), .ZN(n_0_53_12));
   INV_X1 i_0_53_25 (.A(n_0_53_12), .ZN(n_0_1285));
   AOI222_X1 i_0_53_26 (.A1(n_0_1272), .A2(n_0_1252), .B1(n_0_1273), .B2(
      n_0_1220), .C1(n_0_1271), .C2(n_0_1189), .ZN(n_0_53_13));
   INV_X1 i_0_53_27 (.A(n_0_53_13), .ZN(n_0_1286));
   AOI222_X1 i_0_53_28 (.A1(n_0_1272), .A2(n_0_1253), .B1(n_0_1273), .B2(
      n_0_1221), .C1(n_0_1271), .C2(n_0_1190), .ZN(n_0_53_14));
   INV_X1 i_0_53_29 (.A(n_0_53_14), .ZN(n_0_1287));
   AOI222_X1 i_0_53_30 (.A1(n_0_1272), .A2(n_0_1254), .B1(n_0_1273), .B2(
      n_0_1222), .C1(n_0_1271), .C2(n_0_1191), .ZN(n_0_53_15));
   INV_X1 i_0_53_31 (.A(n_0_53_15), .ZN(n_0_1288));
   AOI222_X1 i_0_53_32 (.A1(n_0_1272), .A2(n_0_1255), .B1(n_0_1273), .B2(
      n_0_1223), .C1(n_0_1271), .C2(n_0_1192), .ZN(n_0_53_16));
   INV_X1 i_0_53_33 (.A(n_0_53_16), .ZN(n_0_1289));
   AOI222_X1 i_0_53_34 (.A1(n_0_1272), .A2(n_0_1256), .B1(n_0_1273), .B2(
      n_0_1224), .C1(n_0_1271), .C2(n_0_1193), .ZN(n_0_53_17));
   INV_X1 i_0_53_35 (.A(n_0_53_17), .ZN(n_0_1290));
   AOI222_X1 i_0_53_36 (.A1(n_0_1272), .A2(n_0_1257), .B1(n_0_1273), .B2(
      n_0_1225), .C1(n_0_1271), .C2(n_0_1194), .ZN(n_0_53_18));
   INV_X1 i_0_53_37 (.A(n_0_53_18), .ZN(n_0_1291));
   AOI222_X1 i_0_53_38 (.A1(n_0_1272), .A2(n_0_1258), .B1(n_0_1273), .B2(
      n_0_1226), .C1(n_0_1271), .C2(n_0_1195), .ZN(n_0_53_19));
   INV_X1 i_0_53_39 (.A(n_0_53_19), .ZN(n_0_1292));
   AOI222_X1 i_0_53_40 (.A1(n_0_1272), .A2(n_0_1259), .B1(n_0_1273), .B2(
      n_0_1227), .C1(n_0_1271), .C2(n_0_1196), .ZN(n_0_53_20));
   INV_X1 i_0_53_41 (.A(n_0_53_20), .ZN(n_0_1293));
   AOI222_X1 i_0_53_42 (.A1(n_0_1272), .A2(n_0_1260), .B1(n_0_1273), .B2(
      n_0_1228), .C1(n_0_1271), .C2(n_0_1197), .ZN(n_0_53_21));
   INV_X1 i_0_53_43 (.A(n_0_53_21), .ZN(n_0_1294));
   AOI222_X1 i_0_53_44 (.A1(n_0_1272), .A2(n_0_1261), .B1(n_0_1273), .B2(
      n_0_1229), .C1(n_0_1271), .C2(n_0_1198), .ZN(n_0_53_22));
   INV_X1 i_0_53_45 (.A(n_0_53_22), .ZN(n_0_1295));
   AOI222_X1 i_0_53_46 (.A1(n_0_1272), .A2(n_0_1262), .B1(n_0_1273), .B2(
      n_0_1230), .C1(n_0_1271), .C2(n_0_1199), .ZN(n_0_53_23));
   INV_X1 i_0_53_47 (.A(n_0_53_23), .ZN(n_0_1296));
   AOI222_X1 i_0_53_48 (.A1(n_0_1272), .A2(n_0_1263), .B1(n_0_1273), .B2(
      n_0_1231), .C1(n_0_1271), .C2(n_0_1200), .ZN(n_0_53_24));
   INV_X1 i_0_53_49 (.A(n_0_53_24), .ZN(n_0_1297));
   AOI222_X1 i_0_53_50 (.A1(n_0_1272), .A2(n_0_1264), .B1(n_0_1273), .B2(
      n_0_1232), .C1(n_0_1271), .C2(n_0_1201), .ZN(n_0_53_25));
   INV_X1 i_0_53_51 (.A(n_0_53_25), .ZN(n_0_1298));
   AOI222_X1 i_0_53_52 (.A1(n_0_1272), .A2(n_0_1265), .B1(n_0_1273), .B2(
      n_0_1233), .C1(n_0_1271), .C2(n_0_1202), .ZN(n_0_53_26));
   INV_X1 i_0_53_53 (.A(n_0_53_26), .ZN(n_0_1299));
   AOI222_X1 i_0_53_54 (.A1(n_0_1272), .A2(n_0_1266), .B1(n_0_1273), .B2(
      n_0_1234), .C1(n_0_1271), .C2(n_0_1203), .ZN(n_0_53_27));
   INV_X1 i_0_53_55 (.A(n_0_53_27), .ZN(n_0_1300));
   AOI222_X1 i_0_53_56 (.A1(n_0_1272), .A2(n_0_1267), .B1(n_0_1273), .B2(
      n_0_1235), .C1(n_0_1271), .C2(n_0_1204), .ZN(n_0_53_28));
   INV_X1 i_0_53_57 (.A(n_0_53_28), .ZN(n_0_1301));
   AOI222_X1 i_0_53_58 (.A1(n_0_1272), .A2(n_0_1268), .B1(n_0_1273), .B2(
      n_0_1236), .C1(n_0_1271), .C2(n_0_1205), .ZN(n_0_53_29));
   INV_X1 i_0_53_59 (.A(n_0_53_29), .ZN(n_0_1302));
   AND2_X1 i_0_53_60 (.A1(n_0_1271), .A2(n_0_1206), .ZN(n_0_53_30));
   AOI221_X1 i_0_53_61 (.A(n_0_53_30), .B1(n_0_1272), .B2(n_0_1269), .C1(
      n_0_1273), .C2(n_0_1237), .ZN(n_0_53_31));
   INV_X1 i_0_53_62 (.A(n_0_53_31), .ZN(n_0_1303));
   AOI221_X1 i_0_53_63 (.A(n_0_53_30), .B1(n_0_1272), .B2(n_0_1270), .C1(
      n_0_1273), .C2(n_0_1238), .ZN(n_0_53_32));
   INV_X1 i_0_53_64 (.A(n_0_53_32), .ZN(n_0_1304));
   datapath__0_52 i_0_54 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_27, 
      n_0_1304, n_0_1303, n_0_1302, n_0_1301, n_0_1300, n_0_1299, n_0_1298, 
      n_0_1297, n_0_1296, n_0_1295, n_0_1294, n_0_1293, n_0_1292, n_0_1291, 
      n_0_1290, n_0_1289, n_0_1288, n_0_1287, n_0_1286, n_0_1285, n_0_1284, 
      n_0_1283, n_0_1282, n_0_1281, n_0_1280, n_0_1279, n_0_1278, n_0_1277, 
      n_0_1276, n_0_1275, n_0_1274}), .p_2({n_0_1336, n_0_1335, n_0_1334, 
      n_0_1333, n_0_1332, n_0_1331, n_0_1330, n_0_1329, n_0_1328, n_0_1327, 
      n_0_1326, n_0_1325, n_0_1324, n_0_1323, n_0_1322, n_0_1321, n_0_1320, 
      n_0_1319, n_0_1318, n_0_1317, n_0_1316, n_0_1315, n_0_1314, n_0_1313, 
      n_0_1312, n_0_1311, n_0_1310, n_0_1309, n_0_1308, n_0_1307, n_0_1306, 
      n_0_1305}));
   datapath__0_53 i_0_55 (.multiplicand2(multiplicand2), .p_0({uc_28, n_0_1304, 
      n_0_1303, n_0_1302, n_0_1301, n_0_1300, n_0_1299, n_0_1298, n_0_1297, 
      n_0_1296, n_0_1295, n_0_1294, n_0_1293, n_0_1292, n_0_1291, n_0_1290, 
      n_0_1289, n_0_1288, n_0_1287, n_0_1286, n_0_1285, n_0_1284, n_0_1283, 
      n_0_1282, n_0_1281, n_0_1280, n_0_1279, n_0_1278, n_0_1277, n_0_1276, 
      n_0_1275, n_0_1274}), .p_1({n_0_1368, n_0_1367, n_0_1366, n_0_1365, 
      n_0_1364, n_0_1363, n_0_1362, n_0_1361, n_0_1360, n_0_1359, n_0_1358, 
      n_0_1357, n_0_1356, n_0_1355, n_0_1354, n_0_1353, n_0_1352, n_0_1351, 
      n_0_1350, n_0_1349, n_0_1348, n_0_1347, n_0_1346, n_0_1345, n_0_1344, 
      n_0_1343, n_0_1342, n_0_1341, n_0_1340, n_0_1339, n_0_1338, n_0_1337}));
   INV_X1 i_0_56_0 (.A(multiplier2[14]), .ZN(n_0_56_0));
   AND2_X1 i_0_56_1 (.A1(n_0_56_0), .A2(multiplier2[13]), .ZN(n_0_1370));
   NOR2_X1 i_0_56_2 (.A1(n_0_56_0), .A2(multiplier2[13]), .ZN(n_0_1371));
   NOR2_X1 i_0_56_3 (.A1(n_0_1370), .A2(n_0_1371), .ZN(n_0_1369));
   AOI222_X1 i_0_57_0 (.A1(n_0_1337), .A2(n_0_1370), .B1(n_0_1305), .B2(n_0_1371), 
      .C1(n_0_1274), .C2(n_0_1369), .ZN(n_0_57_0));
   INV_X1 i_0_57_1 (.A(n_0_57_0), .ZN(product[14]));
   AOI222_X1 i_0_57_2 (.A1(n_0_1370), .A2(n_0_1338), .B1(n_0_1371), .B2(n_0_1306), 
      .C1(n_0_1369), .C2(n_0_1275), .ZN(n_0_57_1));
   INV_X1 i_0_57_3 (.A(n_0_57_1), .ZN(n_0_1372));
   AOI222_X1 i_0_57_4 (.A1(n_0_1370), .A2(n_0_1339), .B1(n_0_1371), .B2(n_0_1307), 
      .C1(n_0_1369), .C2(n_0_1276), .ZN(n_0_57_2));
   INV_X1 i_0_57_5 (.A(n_0_57_2), .ZN(n_0_1373));
   AOI222_X1 i_0_57_6 (.A1(n_0_1370), .A2(n_0_1340), .B1(n_0_1371), .B2(n_0_1308), 
      .C1(n_0_1369), .C2(n_0_1277), .ZN(n_0_57_3));
   INV_X1 i_0_57_7 (.A(n_0_57_3), .ZN(n_0_1374));
   AOI222_X1 i_0_57_8 (.A1(n_0_1370), .A2(n_0_1341), .B1(n_0_1371), .B2(n_0_1309), 
      .C1(n_0_1369), .C2(n_0_1278), .ZN(n_0_57_4));
   INV_X1 i_0_57_9 (.A(n_0_57_4), .ZN(n_0_1375));
   AOI222_X1 i_0_57_10 (.A1(n_0_1370), .A2(n_0_1342), .B1(n_0_1371), .B2(
      n_0_1310), .C1(n_0_1369), .C2(n_0_1279), .ZN(n_0_57_5));
   INV_X1 i_0_57_11 (.A(n_0_57_5), .ZN(n_0_1376));
   AOI222_X1 i_0_57_12 (.A1(n_0_1370), .A2(n_0_1343), .B1(n_0_1371), .B2(
      n_0_1311), .C1(n_0_1369), .C2(n_0_1280), .ZN(n_0_57_6));
   INV_X1 i_0_57_13 (.A(n_0_57_6), .ZN(n_0_1377));
   AOI222_X1 i_0_57_14 (.A1(n_0_1370), .A2(n_0_1344), .B1(n_0_1371), .B2(
      n_0_1312), .C1(n_0_1369), .C2(n_0_1281), .ZN(n_0_57_7));
   INV_X1 i_0_57_15 (.A(n_0_57_7), .ZN(n_0_1378));
   AOI222_X1 i_0_57_16 (.A1(n_0_1370), .A2(n_0_1345), .B1(n_0_1371), .B2(
      n_0_1313), .C1(n_0_1369), .C2(n_0_1282), .ZN(n_0_57_8));
   INV_X1 i_0_57_17 (.A(n_0_57_8), .ZN(n_0_1379));
   AOI222_X1 i_0_57_18 (.A1(n_0_1370), .A2(n_0_1346), .B1(n_0_1371), .B2(
      n_0_1314), .C1(n_0_1369), .C2(n_0_1283), .ZN(n_0_57_9));
   INV_X1 i_0_57_19 (.A(n_0_57_9), .ZN(n_0_1380));
   AOI222_X1 i_0_57_20 (.A1(n_0_1370), .A2(n_0_1347), .B1(n_0_1371), .B2(
      n_0_1315), .C1(n_0_1369), .C2(n_0_1284), .ZN(n_0_57_10));
   INV_X1 i_0_57_21 (.A(n_0_57_10), .ZN(n_0_1381));
   AOI222_X1 i_0_57_22 (.A1(n_0_1370), .A2(n_0_1348), .B1(n_0_1371), .B2(
      n_0_1316), .C1(n_0_1369), .C2(n_0_1285), .ZN(n_0_57_11));
   INV_X1 i_0_57_23 (.A(n_0_57_11), .ZN(n_0_1382));
   AOI222_X1 i_0_57_24 (.A1(n_0_1370), .A2(n_0_1349), .B1(n_0_1371), .B2(
      n_0_1317), .C1(n_0_1369), .C2(n_0_1286), .ZN(n_0_57_12));
   INV_X1 i_0_57_25 (.A(n_0_57_12), .ZN(n_0_1383));
   AOI222_X1 i_0_57_26 (.A1(n_0_1370), .A2(n_0_1350), .B1(n_0_1371), .B2(
      n_0_1318), .C1(n_0_1369), .C2(n_0_1287), .ZN(n_0_57_13));
   INV_X1 i_0_57_27 (.A(n_0_57_13), .ZN(n_0_1384));
   AOI222_X1 i_0_57_28 (.A1(n_0_1370), .A2(n_0_1351), .B1(n_0_1371), .B2(
      n_0_1319), .C1(n_0_1369), .C2(n_0_1288), .ZN(n_0_57_14));
   INV_X1 i_0_57_29 (.A(n_0_57_14), .ZN(n_0_1385));
   AOI222_X1 i_0_57_30 (.A1(n_0_1370), .A2(n_0_1352), .B1(n_0_1371), .B2(
      n_0_1320), .C1(n_0_1369), .C2(n_0_1289), .ZN(n_0_57_15));
   INV_X1 i_0_57_31 (.A(n_0_57_15), .ZN(n_0_1386));
   AOI222_X1 i_0_57_32 (.A1(n_0_1370), .A2(n_0_1353), .B1(n_0_1371), .B2(
      n_0_1321), .C1(n_0_1369), .C2(n_0_1290), .ZN(n_0_57_16));
   INV_X1 i_0_57_33 (.A(n_0_57_16), .ZN(n_0_1387));
   AOI222_X1 i_0_57_34 (.A1(n_0_1370), .A2(n_0_1354), .B1(n_0_1371), .B2(
      n_0_1322), .C1(n_0_1369), .C2(n_0_1291), .ZN(n_0_57_17));
   INV_X1 i_0_57_35 (.A(n_0_57_17), .ZN(n_0_1388));
   AOI222_X1 i_0_57_36 (.A1(n_0_1370), .A2(n_0_1355), .B1(n_0_1371), .B2(
      n_0_1323), .C1(n_0_1369), .C2(n_0_1292), .ZN(n_0_57_18));
   INV_X1 i_0_57_37 (.A(n_0_57_18), .ZN(n_0_1389));
   AOI222_X1 i_0_57_38 (.A1(n_0_1370), .A2(n_0_1356), .B1(n_0_1371), .B2(
      n_0_1324), .C1(n_0_1369), .C2(n_0_1293), .ZN(n_0_57_19));
   INV_X1 i_0_57_39 (.A(n_0_57_19), .ZN(n_0_1390));
   AOI222_X1 i_0_57_40 (.A1(n_0_1370), .A2(n_0_1357), .B1(n_0_1371), .B2(
      n_0_1325), .C1(n_0_1369), .C2(n_0_1294), .ZN(n_0_57_20));
   INV_X1 i_0_57_41 (.A(n_0_57_20), .ZN(n_0_1391));
   AOI222_X1 i_0_57_42 (.A1(n_0_1370), .A2(n_0_1358), .B1(n_0_1371), .B2(
      n_0_1326), .C1(n_0_1369), .C2(n_0_1295), .ZN(n_0_57_21));
   INV_X1 i_0_57_43 (.A(n_0_57_21), .ZN(n_0_1392));
   AOI222_X1 i_0_57_44 (.A1(n_0_1370), .A2(n_0_1359), .B1(n_0_1371), .B2(
      n_0_1327), .C1(n_0_1369), .C2(n_0_1296), .ZN(n_0_57_22));
   INV_X1 i_0_57_45 (.A(n_0_57_22), .ZN(n_0_1393));
   AOI222_X1 i_0_57_46 (.A1(n_0_1370), .A2(n_0_1360), .B1(n_0_1371), .B2(
      n_0_1328), .C1(n_0_1369), .C2(n_0_1297), .ZN(n_0_57_23));
   INV_X1 i_0_57_47 (.A(n_0_57_23), .ZN(n_0_1394));
   AOI222_X1 i_0_57_48 (.A1(n_0_1370), .A2(n_0_1361), .B1(n_0_1371), .B2(
      n_0_1329), .C1(n_0_1369), .C2(n_0_1298), .ZN(n_0_57_24));
   INV_X1 i_0_57_49 (.A(n_0_57_24), .ZN(n_0_1395));
   AOI222_X1 i_0_57_50 (.A1(n_0_1370), .A2(n_0_1362), .B1(n_0_1371), .B2(
      n_0_1330), .C1(n_0_1369), .C2(n_0_1299), .ZN(n_0_57_25));
   INV_X1 i_0_57_51 (.A(n_0_57_25), .ZN(n_0_1396));
   AOI222_X1 i_0_57_52 (.A1(n_0_1370), .A2(n_0_1363), .B1(n_0_1371), .B2(
      n_0_1331), .C1(n_0_1369), .C2(n_0_1300), .ZN(n_0_57_26));
   INV_X1 i_0_57_53 (.A(n_0_57_26), .ZN(n_0_1397));
   AOI222_X1 i_0_57_54 (.A1(n_0_1370), .A2(n_0_1364), .B1(n_0_1371), .B2(
      n_0_1332), .C1(n_0_1369), .C2(n_0_1301), .ZN(n_0_57_27));
   INV_X1 i_0_57_55 (.A(n_0_57_27), .ZN(n_0_1398));
   AOI222_X1 i_0_57_56 (.A1(n_0_1370), .A2(n_0_1365), .B1(n_0_1371), .B2(
      n_0_1333), .C1(n_0_1369), .C2(n_0_1302), .ZN(n_0_57_28));
   INV_X1 i_0_57_57 (.A(n_0_57_28), .ZN(n_0_1399));
   AOI222_X1 i_0_57_58 (.A1(n_0_1370), .A2(n_0_1366), .B1(n_0_1371), .B2(
      n_0_1334), .C1(n_0_1369), .C2(n_0_1303), .ZN(n_0_57_29));
   INV_X1 i_0_57_59 (.A(n_0_57_29), .ZN(n_0_1400));
   AND2_X1 i_0_57_60 (.A1(n_0_1369), .A2(n_0_1304), .ZN(n_0_57_30));
   AOI221_X1 i_0_57_61 (.A(n_0_57_30), .B1(n_0_1370), .B2(n_0_1367), .C1(
      n_0_1371), .C2(n_0_1335), .ZN(n_0_57_31));
   INV_X1 i_0_57_62 (.A(n_0_57_31), .ZN(n_0_1401));
   AOI221_X1 i_0_57_63 (.A(n_0_57_30), .B1(n_0_1370), .B2(n_0_1368), .C1(
      n_0_1371), .C2(n_0_1336), .ZN(n_0_57_32));
   INV_X1 i_0_57_64 (.A(n_0_57_32), .ZN(n_0_1402));
   datapath__0_56 i_0_58 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_29, 
      n_0_1402, n_0_1401, n_0_1400, n_0_1399, n_0_1398, n_0_1397, n_0_1396, 
      n_0_1395, n_0_1394, n_0_1393, n_0_1392, n_0_1391, n_0_1390, n_0_1389, 
      n_0_1388, n_0_1387, n_0_1386, n_0_1385, n_0_1384, n_0_1383, n_0_1382, 
      n_0_1381, n_0_1380, n_0_1379, n_0_1378, n_0_1377, n_0_1376, n_0_1375, 
      n_0_1374, n_0_1373, n_0_1372}), .p_2({n_0_1434, n_0_1433, n_0_1432, 
      n_0_1431, n_0_1430, n_0_1429, n_0_1428, n_0_1427, n_0_1426, n_0_1425, 
      n_0_1424, n_0_1423, n_0_1422, n_0_1421, n_0_1420, n_0_1419, n_0_1418, 
      n_0_1417, n_0_1416, n_0_1415, n_0_1414, n_0_1413, n_0_1412, n_0_1411, 
      n_0_1410, n_0_1409, n_0_1408, n_0_1407, n_0_1406, n_0_1405, n_0_1404, 
      n_0_1403}));
   datapath__0_57 i_0_59 (.multiplicand2(multiplicand2), .p_0({uc_30, n_0_1402, 
      n_0_1401, n_0_1400, n_0_1399, n_0_1398, n_0_1397, n_0_1396, n_0_1395, 
      n_0_1394, n_0_1393, n_0_1392, n_0_1391, n_0_1390, n_0_1389, n_0_1388, 
      n_0_1387, n_0_1386, n_0_1385, n_0_1384, n_0_1383, n_0_1382, n_0_1381, 
      n_0_1380, n_0_1379, n_0_1378, n_0_1377, n_0_1376, n_0_1375, n_0_1374, 
      n_0_1373, n_0_1372}), .p_1({n_0_1466, n_0_1465, n_0_1464, n_0_1463, 
      n_0_1462, n_0_1461, n_0_1460, n_0_1459, n_0_1458, n_0_1457, n_0_1456, 
      n_0_1455, n_0_1454, n_0_1453, n_0_1452, n_0_1451, n_0_1450, n_0_1449, 
      n_0_1448, n_0_1447, n_0_1446, n_0_1445, n_0_1444, n_0_1443, n_0_1442, 
      n_0_1441, n_0_1440, n_0_1439, n_0_1438, n_0_1437, n_0_1436, n_0_1435}));
   INV_X1 i_0_60_0 (.A(multiplier2[15]), .ZN(n_0_60_0));
   AND2_X1 i_0_60_1 (.A1(n_0_60_0), .A2(multiplier2[14]), .ZN(n_0_1468));
   NOR2_X1 i_0_60_2 (.A1(n_0_60_0), .A2(multiplier2[14]), .ZN(n_0_1469));
   NOR2_X1 i_0_60_3 (.A1(n_0_1468), .A2(n_0_1469), .ZN(n_0_1467));
   AOI222_X1 i_0_61_0 (.A1(n_0_1435), .A2(n_0_1468), .B1(n_0_1403), .B2(n_0_1469), 
      .C1(n_0_1372), .C2(n_0_1467), .ZN(n_0_61_0));
   INV_X1 i_0_61_1 (.A(n_0_61_0), .ZN(product[15]));
   AOI222_X1 i_0_61_2 (.A1(n_0_1468), .A2(n_0_1436), .B1(n_0_1469), .B2(n_0_1404), 
      .C1(n_0_1467), .C2(n_0_1373), .ZN(n_0_61_1));
   INV_X1 i_0_61_3 (.A(n_0_61_1), .ZN(n_0_1470));
   AOI222_X1 i_0_61_4 (.A1(n_0_1468), .A2(n_0_1437), .B1(n_0_1469), .B2(n_0_1405), 
      .C1(n_0_1467), .C2(n_0_1374), .ZN(n_0_61_2));
   INV_X1 i_0_61_5 (.A(n_0_61_2), .ZN(n_0_1471));
   AOI222_X1 i_0_61_6 (.A1(n_0_1468), .A2(n_0_1438), .B1(n_0_1469), .B2(n_0_1406), 
      .C1(n_0_1467), .C2(n_0_1375), .ZN(n_0_61_3));
   INV_X1 i_0_61_7 (.A(n_0_61_3), .ZN(n_0_1472));
   AOI222_X1 i_0_61_8 (.A1(n_0_1468), .A2(n_0_1439), .B1(n_0_1469), .B2(n_0_1407), 
      .C1(n_0_1467), .C2(n_0_1376), .ZN(n_0_61_4));
   INV_X1 i_0_61_9 (.A(n_0_61_4), .ZN(n_0_1473));
   AOI222_X1 i_0_61_10 (.A1(n_0_1468), .A2(n_0_1440), .B1(n_0_1469), .B2(
      n_0_1408), .C1(n_0_1467), .C2(n_0_1377), .ZN(n_0_61_5));
   INV_X1 i_0_61_11 (.A(n_0_61_5), .ZN(n_0_1474));
   AOI222_X1 i_0_61_12 (.A1(n_0_1468), .A2(n_0_1441), .B1(n_0_1469), .B2(
      n_0_1409), .C1(n_0_1467), .C2(n_0_1378), .ZN(n_0_61_6));
   INV_X1 i_0_61_13 (.A(n_0_61_6), .ZN(n_0_1475));
   AOI222_X1 i_0_61_14 (.A1(n_0_1468), .A2(n_0_1442), .B1(n_0_1469), .B2(
      n_0_1410), .C1(n_0_1467), .C2(n_0_1379), .ZN(n_0_61_7));
   INV_X1 i_0_61_15 (.A(n_0_61_7), .ZN(n_0_1476));
   AOI222_X1 i_0_61_16 (.A1(n_0_1468), .A2(n_0_1443), .B1(n_0_1469), .B2(
      n_0_1411), .C1(n_0_1467), .C2(n_0_1380), .ZN(n_0_61_8));
   INV_X1 i_0_61_17 (.A(n_0_61_8), .ZN(n_0_1477));
   AOI222_X1 i_0_61_18 (.A1(n_0_1468), .A2(n_0_1444), .B1(n_0_1469), .B2(
      n_0_1412), .C1(n_0_1467), .C2(n_0_1381), .ZN(n_0_61_9));
   INV_X1 i_0_61_19 (.A(n_0_61_9), .ZN(n_0_1478));
   AOI222_X1 i_0_61_20 (.A1(n_0_1468), .A2(n_0_1445), .B1(n_0_1469), .B2(
      n_0_1413), .C1(n_0_1467), .C2(n_0_1382), .ZN(n_0_61_10));
   INV_X1 i_0_61_21 (.A(n_0_61_10), .ZN(n_0_1479));
   AOI222_X1 i_0_61_22 (.A1(n_0_1468), .A2(n_0_1446), .B1(n_0_1469), .B2(
      n_0_1414), .C1(n_0_1467), .C2(n_0_1383), .ZN(n_0_61_11));
   INV_X1 i_0_61_23 (.A(n_0_61_11), .ZN(n_0_1480));
   AOI222_X1 i_0_61_24 (.A1(n_0_1468), .A2(n_0_1447), .B1(n_0_1469), .B2(
      n_0_1415), .C1(n_0_1467), .C2(n_0_1384), .ZN(n_0_61_12));
   INV_X1 i_0_61_25 (.A(n_0_61_12), .ZN(n_0_1481));
   AOI222_X1 i_0_61_26 (.A1(n_0_1468), .A2(n_0_1448), .B1(n_0_1469), .B2(
      n_0_1416), .C1(n_0_1467), .C2(n_0_1385), .ZN(n_0_61_13));
   INV_X1 i_0_61_27 (.A(n_0_61_13), .ZN(n_0_1482));
   AOI222_X1 i_0_61_28 (.A1(n_0_1468), .A2(n_0_1449), .B1(n_0_1469), .B2(
      n_0_1417), .C1(n_0_1467), .C2(n_0_1386), .ZN(n_0_61_14));
   INV_X1 i_0_61_29 (.A(n_0_61_14), .ZN(n_0_1483));
   AOI222_X1 i_0_61_30 (.A1(n_0_1468), .A2(n_0_1450), .B1(n_0_1469), .B2(
      n_0_1418), .C1(n_0_1467), .C2(n_0_1387), .ZN(n_0_61_15));
   INV_X1 i_0_61_31 (.A(n_0_61_15), .ZN(n_0_1484));
   AOI222_X1 i_0_61_32 (.A1(n_0_1468), .A2(n_0_1451), .B1(n_0_1469), .B2(
      n_0_1419), .C1(n_0_1467), .C2(n_0_1388), .ZN(n_0_61_16));
   INV_X1 i_0_61_33 (.A(n_0_61_16), .ZN(n_0_1485));
   AOI222_X1 i_0_61_34 (.A1(n_0_1468), .A2(n_0_1452), .B1(n_0_1469), .B2(
      n_0_1420), .C1(n_0_1467), .C2(n_0_1389), .ZN(n_0_61_17));
   INV_X1 i_0_61_35 (.A(n_0_61_17), .ZN(n_0_1486));
   AOI222_X1 i_0_61_36 (.A1(n_0_1468), .A2(n_0_1453), .B1(n_0_1469), .B2(
      n_0_1421), .C1(n_0_1467), .C2(n_0_1390), .ZN(n_0_61_18));
   INV_X1 i_0_61_37 (.A(n_0_61_18), .ZN(n_0_1487));
   AOI222_X1 i_0_61_38 (.A1(n_0_1468), .A2(n_0_1454), .B1(n_0_1469), .B2(
      n_0_1422), .C1(n_0_1467), .C2(n_0_1391), .ZN(n_0_61_19));
   INV_X1 i_0_61_39 (.A(n_0_61_19), .ZN(n_0_1488));
   AOI222_X1 i_0_61_40 (.A1(n_0_1468), .A2(n_0_1455), .B1(n_0_1469), .B2(
      n_0_1423), .C1(n_0_1467), .C2(n_0_1392), .ZN(n_0_61_20));
   INV_X1 i_0_61_41 (.A(n_0_61_20), .ZN(n_0_1489));
   AOI222_X1 i_0_61_42 (.A1(n_0_1468), .A2(n_0_1456), .B1(n_0_1469), .B2(
      n_0_1424), .C1(n_0_1467), .C2(n_0_1393), .ZN(n_0_61_21));
   INV_X1 i_0_61_43 (.A(n_0_61_21), .ZN(n_0_1490));
   AOI222_X1 i_0_61_44 (.A1(n_0_1468), .A2(n_0_1457), .B1(n_0_1469), .B2(
      n_0_1425), .C1(n_0_1467), .C2(n_0_1394), .ZN(n_0_61_22));
   INV_X1 i_0_61_45 (.A(n_0_61_22), .ZN(n_0_1491));
   AOI222_X1 i_0_61_46 (.A1(n_0_1468), .A2(n_0_1458), .B1(n_0_1469), .B2(
      n_0_1426), .C1(n_0_1467), .C2(n_0_1395), .ZN(n_0_61_23));
   INV_X1 i_0_61_47 (.A(n_0_61_23), .ZN(n_0_1492));
   AOI222_X1 i_0_61_48 (.A1(n_0_1468), .A2(n_0_1459), .B1(n_0_1469), .B2(
      n_0_1427), .C1(n_0_1467), .C2(n_0_1396), .ZN(n_0_61_24));
   INV_X1 i_0_61_49 (.A(n_0_61_24), .ZN(n_0_1493));
   AOI222_X1 i_0_61_50 (.A1(n_0_1468), .A2(n_0_1460), .B1(n_0_1469), .B2(
      n_0_1428), .C1(n_0_1467), .C2(n_0_1397), .ZN(n_0_61_25));
   INV_X1 i_0_61_51 (.A(n_0_61_25), .ZN(n_0_1494));
   AOI222_X1 i_0_61_52 (.A1(n_0_1468), .A2(n_0_1461), .B1(n_0_1469), .B2(
      n_0_1429), .C1(n_0_1467), .C2(n_0_1398), .ZN(n_0_61_26));
   INV_X1 i_0_61_53 (.A(n_0_61_26), .ZN(n_0_1495));
   AOI222_X1 i_0_61_54 (.A1(n_0_1468), .A2(n_0_1462), .B1(n_0_1469), .B2(
      n_0_1430), .C1(n_0_1467), .C2(n_0_1399), .ZN(n_0_61_27));
   INV_X1 i_0_61_55 (.A(n_0_61_27), .ZN(n_0_1496));
   AOI222_X1 i_0_61_56 (.A1(n_0_1468), .A2(n_0_1463), .B1(n_0_1469), .B2(
      n_0_1431), .C1(n_0_1467), .C2(n_0_1400), .ZN(n_0_61_28));
   INV_X1 i_0_61_57 (.A(n_0_61_28), .ZN(n_0_1497));
   AOI222_X1 i_0_61_58 (.A1(n_0_1468), .A2(n_0_1464), .B1(n_0_1469), .B2(
      n_0_1432), .C1(n_0_1467), .C2(n_0_1401), .ZN(n_0_61_29));
   INV_X1 i_0_61_59 (.A(n_0_61_29), .ZN(n_0_1498));
   AND2_X1 i_0_61_60 (.A1(n_0_1467), .A2(n_0_1402), .ZN(n_0_61_30));
   AOI221_X1 i_0_61_61 (.A(n_0_61_30), .B1(n_0_1468), .B2(n_0_1465), .C1(
      n_0_1469), .C2(n_0_1433), .ZN(n_0_61_31));
   INV_X1 i_0_61_62 (.A(n_0_61_31), .ZN(n_0_1499));
   AOI221_X1 i_0_61_63 (.A(n_0_61_30), .B1(n_0_1468), .B2(n_0_1466), .C1(
      n_0_1469), .C2(n_0_1434), .ZN(n_0_61_32));
   INV_X1 i_0_61_64 (.A(n_0_61_32), .ZN(n_0_1500));
   datapath__0_60 i_0_62 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_31, 
      n_0_1500, n_0_1499, n_0_1498, n_0_1497, n_0_1496, n_0_1495, n_0_1494, 
      n_0_1493, n_0_1492, n_0_1491, n_0_1490, n_0_1489, n_0_1488, n_0_1487, 
      n_0_1486, n_0_1485, n_0_1484, n_0_1483, n_0_1482, n_0_1481, n_0_1480, 
      n_0_1479, n_0_1478, n_0_1477, n_0_1476, n_0_1475, n_0_1474, n_0_1473, 
      n_0_1472, n_0_1471, n_0_1470}), .p_2({n_0_1532, n_0_1531, n_0_1530, 
      n_0_1529, n_0_1528, n_0_1527, n_0_1526, n_0_1525, n_0_1524, n_0_1523, 
      n_0_1522, n_0_1521, n_0_1520, n_0_1519, n_0_1518, n_0_1517, n_0_1516, 
      n_0_1515, n_0_1514, n_0_1513, n_0_1512, n_0_1511, n_0_1510, n_0_1509, 
      n_0_1508, n_0_1507, n_0_1506, n_0_1505, n_0_1504, n_0_1503, n_0_1502, 
      n_0_1501}));
   datapath__0_61 i_0_63 (.multiplicand2(multiplicand2), .p_0({uc_32, n_0_1500, 
      n_0_1499, n_0_1498, n_0_1497, n_0_1496, n_0_1495, n_0_1494, n_0_1493, 
      n_0_1492, n_0_1491, n_0_1490, n_0_1489, n_0_1488, n_0_1487, n_0_1486, 
      n_0_1485, n_0_1484, n_0_1483, n_0_1482, n_0_1481, n_0_1480, n_0_1479, 
      n_0_1478, n_0_1477, n_0_1476, n_0_1475, n_0_1474, n_0_1473, n_0_1472, 
      n_0_1471, n_0_1470}), .p_1({n_0_1564, n_0_1563, n_0_1562, n_0_1561, 
      n_0_1560, n_0_1559, n_0_1558, n_0_1557, n_0_1556, n_0_1555, n_0_1554, 
      n_0_1553, n_0_1552, n_0_1551, n_0_1550, n_0_1549, n_0_1548, n_0_1547, 
      n_0_1546, n_0_1545, n_0_1544, n_0_1543, n_0_1542, n_0_1541, n_0_1540, 
      n_0_1539, n_0_1538, n_0_1537, n_0_1536, n_0_1535, n_0_1534, n_0_1533}));
   INV_X1 i_0_64_0 (.A(multiplier2[16]), .ZN(n_0_64_0));
   AND2_X1 i_0_64_1 (.A1(n_0_64_0), .A2(multiplier2[15]), .ZN(n_0_1566));
   NOR2_X1 i_0_64_2 (.A1(n_0_64_0), .A2(multiplier2[15]), .ZN(n_0_1567));
   NOR2_X1 i_0_64_3 (.A1(n_0_1566), .A2(n_0_1567), .ZN(n_0_1565));
   AOI222_X1 i_0_65_0 (.A1(n_0_1533), .A2(n_0_1566), .B1(n_0_1501), .B2(n_0_1567), 
      .C1(n_0_1470), .C2(n_0_1565), .ZN(n_0_65_0));
   INV_X1 i_0_65_1 (.A(n_0_65_0), .ZN(product[16]));
   AOI222_X1 i_0_65_2 (.A1(n_0_1566), .A2(n_0_1534), .B1(n_0_1567), .B2(n_0_1502), 
      .C1(n_0_1565), .C2(n_0_1471), .ZN(n_0_65_1));
   INV_X1 i_0_65_3 (.A(n_0_65_1), .ZN(n_0_1568));
   AOI222_X1 i_0_65_4 (.A1(n_0_1566), .A2(n_0_1535), .B1(n_0_1567), .B2(n_0_1503), 
      .C1(n_0_1565), .C2(n_0_1472), .ZN(n_0_65_2));
   INV_X1 i_0_65_5 (.A(n_0_65_2), .ZN(n_0_1569));
   AOI222_X1 i_0_65_6 (.A1(n_0_1566), .A2(n_0_1536), .B1(n_0_1567), .B2(n_0_1504), 
      .C1(n_0_1565), .C2(n_0_1473), .ZN(n_0_65_3));
   INV_X1 i_0_65_7 (.A(n_0_65_3), .ZN(n_0_1570));
   AOI222_X1 i_0_65_8 (.A1(n_0_1566), .A2(n_0_1537), .B1(n_0_1567), .B2(n_0_1505), 
      .C1(n_0_1565), .C2(n_0_1474), .ZN(n_0_65_4));
   INV_X1 i_0_65_9 (.A(n_0_65_4), .ZN(n_0_1571));
   AOI222_X1 i_0_65_10 (.A1(n_0_1566), .A2(n_0_1538), .B1(n_0_1567), .B2(
      n_0_1506), .C1(n_0_1565), .C2(n_0_1475), .ZN(n_0_65_5));
   INV_X1 i_0_65_11 (.A(n_0_65_5), .ZN(n_0_1572));
   AOI222_X1 i_0_65_12 (.A1(n_0_1566), .A2(n_0_1539), .B1(n_0_1567), .B2(
      n_0_1507), .C1(n_0_1565), .C2(n_0_1476), .ZN(n_0_65_6));
   INV_X1 i_0_65_13 (.A(n_0_65_6), .ZN(n_0_1573));
   AOI222_X1 i_0_65_14 (.A1(n_0_1566), .A2(n_0_1540), .B1(n_0_1567), .B2(
      n_0_1508), .C1(n_0_1565), .C2(n_0_1477), .ZN(n_0_65_7));
   INV_X1 i_0_65_15 (.A(n_0_65_7), .ZN(n_0_1574));
   AOI222_X1 i_0_65_16 (.A1(n_0_1566), .A2(n_0_1541), .B1(n_0_1567), .B2(
      n_0_1509), .C1(n_0_1565), .C2(n_0_1478), .ZN(n_0_65_8));
   INV_X1 i_0_65_17 (.A(n_0_65_8), .ZN(n_0_1575));
   AOI222_X1 i_0_65_18 (.A1(n_0_1566), .A2(n_0_1542), .B1(n_0_1567), .B2(
      n_0_1510), .C1(n_0_1565), .C2(n_0_1479), .ZN(n_0_65_9));
   INV_X1 i_0_65_19 (.A(n_0_65_9), .ZN(n_0_1576));
   AOI222_X1 i_0_65_20 (.A1(n_0_1566), .A2(n_0_1543), .B1(n_0_1567), .B2(
      n_0_1511), .C1(n_0_1565), .C2(n_0_1480), .ZN(n_0_65_10));
   INV_X1 i_0_65_21 (.A(n_0_65_10), .ZN(n_0_1577));
   AOI222_X1 i_0_65_22 (.A1(n_0_1566), .A2(n_0_1544), .B1(n_0_1567), .B2(
      n_0_1512), .C1(n_0_1565), .C2(n_0_1481), .ZN(n_0_65_11));
   INV_X1 i_0_65_23 (.A(n_0_65_11), .ZN(n_0_1578));
   AOI222_X1 i_0_65_24 (.A1(n_0_1566), .A2(n_0_1545), .B1(n_0_1567), .B2(
      n_0_1513), .C1(n_0_1565), .C2(n_0_1482), .ZN(n_0_65_12));
   INV_X1 i_0_65_25 (.A(n_0_65_12), .ZN(n_0_1579));
   AOI222_X1 i_0_65_26 (.A1(n_0_1566), .A2(n_0_1546), .B1(n_0_1567), .B2(
      n_0_1514), .C1(n_0_1565), .C2(n_0_1483), .ZN(n_0_65_13));
   INV_X1 i_0_65_27 (.A(n_0_65_13), .ZN(n_0_1580));
   AOI222_X1 i_0_65_28 (.A1(n_0_1566), .A2(n_0_1547), .B1(n_0_1567), .B2(
      n_0_1515), .C1(n_0_1565), .C2(n_0_1484), .ZN(n_0_65_14));
   INV_X1 i_0_65_29 (.A(n_0_65_14), .ZN(n_0_1581));
   AOI222_X1 i_0_65_30 (.A1(n_0_1566), .A2(n_0_1548), .B1(n_0_1567), .B2(
      n_0_1516), .C1(n_0_1565), .C2(n_0_1485), .ZN(n_0_65_15));
   INV_X1 i_0_65_31 (.A(n_0_65_15), .ZN(n_0_1582));
   AOI222_X1 i_0_65_32 (.A1(n_0_1566), .A2(n_0_1549), .B1(n_0_1567), .B2(
      n_0_1517), .C1(n_0_1565), .C2(n_0_1486), .ZN(n_0_65_16));
   INV_X1 i_0_65_33 (.A(n_0_65_16), .ZN(n_0_1583));
   AOI222_X1 i_0_65_34 (.A1(n_0_1566), .A2(n_0_1550), .B1(n_0_1567), .B2(
      n_0_1518), .C1(n_0_1565), .C2(n_0_1487), .ZN(n_0_65_17));
   INV_X1 i_0_65_35 (.A(n_0_65_17), .ZN(n_0_1584));
   AOI222_X1 i_0_65_36 (.A1(n_0_1566), .A2(n_0_1551), .B1(n_0_1567), .B2(
      n_0_1519), .C1(n_0_1565), .C2(n_0_1488), .ZN(n_0_65_18));
   INV_X1 i_0_65_37 (.A(n_0_65_18), .ZN(n_0_1585));
   AOI222_X1 i_0_65_38 (.A1(n_0_1566), .A2(n_0_1552), .B1(n_0_1567), .B2(
      n_0_1520), .C1(n_0_1565), .C2(n_0_1489), .ZN(n_0_65_19));
   INV_X1 i_0_65_39 (.A(n_0_65_19), .ZN(n_0_1586));
   AOI222_X1 i_0_65_40 (.A1(n_0_1566), .A2(n_0_1553), .B1(n_0_1567), .B2(
      n_0_1521), .C1(n_0_1565), .C2(n_0_1490), .ZN(n_0_65_20));
   INV_X1 i_0_65_41 (.A(n_0_65_20), .ZN(n_0_1587));
   AOI222_X1 i_0_65_42 (.A1(n_0_1566), .A2(n_0_1554), .B1(n_0_1567), .B2(
      n_0_1522), .C1(n_0_1565), .C2(n_0_1491), .ZN(n_0_65_21));
   INV_X1 i_0_65_43 (.A(n_0_65_21), .ZN(n_0_1588));
   AOI222_X1 i_0_65_44 (.A1(n_0_1566), .A2(n_0_1555), .B1(n_0_1567), .B2(
      n_0_1523), .C1(n_0_1565), .C2(n_0_1492), .ZN(n_0_65_22));
   INV_X1 i_0_65_45 (.A(n_0_65_22), .ZN(n_0_1589));
   AOI222_X1 i_0_65_46 (.A1(n_0_1566), .A2(n_0_1556), .B1(n_0_1567), .B2(
      n_0_1524), .C1(n_0_1565), .C2(n_0_1493), .ZN(n_0_65_23));
   INV_X1 i_0_65_47 (.A(n_0_65_23), .ZN(n_0_1590));
   AOI222_X1 i_0_65_48 (.A1(n_0_1566), .A2(n_0_1557), .B1(n_0_1567), .B2(
      n_0_1525), .C1(n_0_1565), .C2(n_0_1494), .ZN(n_0_65_24));
   INV_X1 i_0_65_49 (.A(n_0_65_24), .ZN(n_0_1591));
   AOI222_X1 i_0_65_50 (.A1(n_0_1566), .A2(n_0_1558), .B1(n_0_1567), .B2(
      n_0_1526), .C1(n_0_1565), .C2(n_0_1495), .ZN(n_0_65_25));
   INV_X1 i_0_65_51 (.A(n_0_65_25), .ZN(n_0_1592));
   AOI222_X1 i_0_65_52 (.A1(n_0_1566), .A2(n_0_1559), .B1(n_0_1567), .B2(
      n_0_1527), .C1(n_0_1565), .C2(n_0_1496), .ZN(n_0_65_26));
   INV_X1 i_0_65_53 (.A(n_0_65_26), .ZN(n_0_1593));
   AOI222_X1 i_0_65_54 (.A1(n_0_1566), .A2(n_0_1560), .B1(n_0_1567), .B2(
      n_0_1528), .C1(n_0_1565), .C2(n_0_1497), .ZN(n_0_65_27));
   INV_X1 i_0_65_55 (.A(n_0_65_27), .ZN(n_0_1594));
   AOI222_X1 i_0_65_56 (.A1(n_0_1566), .A2(n_0_1561), .B1(n_0_1567), .B2(
      n_0_1529), .C1(n_0_1565), .C2(n_0_1498), .ZN(n_0_65_28));
   INV_X1 i_0_65_57 (.A(n_0_65_28), .ZN(n_0_1595));
   AOI222_X1 i_0_65_58 (.A1(n_0_1566), .A2(n_0_1562), .B1(n_0_1567), .B2(
      n_0_1530), .C1(n_0_1565), .C2(n_0_1499), .ZN(n_0_65_29));
   INV_X1 i_0_65_59 (.A(n_0_65_29), .ZN(n_0_1596));
   AND2_X1 i_0_65_60 (.A1(n_0_1565), .A2(n_0_1500), .ZN(n_0_65_30));
   AOI221_X1 i_0_65_61 (.A(n_0_65_30), .B1(n_0_1566), .B2(n_0_1563), .C1(
      n_0_1567), .C2(n_0_1531), .ZN(n_0_65_31));
   INV_X1 i_0_65_62 (.A(n_0_65_31), .ZN(n_0_1597));
   AOI221_X1 i_0_65_63 (.A(n_0_65_30), .B1(n_0_1566), .B2(n_0_1564), .C1(
      n_0_1567), .C2(n_0_1532), .ZN(n_0_65_32));
   INV_X1 i_0_65_64 (.A(n_0_65_32), .ZN(n_0_1598));
   datapath__0_64 i_0_66 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_33, 
      n_0_1598, n_0_1597, n_0_1596, n_0_1595, n_0_1594, n_0_1593, n_0_1592, 
      n_0_1591, n_0_1590, n_0_1589, n_0_1588, n_0_1587, n_0_1586, n_0_1585, 
      n_0_1584, n_0_1583, n_0_1582, n_0_1581, n_0_1580, n_0_1579, n_0_1578, 
      n_0_1577, n_0_1576, n_0_1575, n_0_1574, n_0_1573, n_0_1572, n_0_1571, 
      n_0_1570, n_0_1569, n_0_1568}), .p_2({n_0_1630, n_0_1629, n_0_1628, 
      n_0_1627, n_0_1626, n_0_1625, n_0_1624, n_0_1623, n_0_1622, n_0_1621, 
      n_0_1620, n_0_1619, n_0_1618, n_0_1617, n_0_1616, n_0_1615, n_0_1614, 
      n_0_1613, n_0_1612, n_0_1611, n_0_1610, n_0_1609, n_0_1608, n_0_1607, 
      n_0_1606, n_0_1605, n_0_1604, n_0_1603, n_0_1602, n_0_1601, n_0_1600, 
      n_0_1599}));
   datapath__0_65 i_0_67 (.multiplicand2(multiplicand2), .p_0({uc_34, n_0_1598, 
      n_0_1597, n_0_1596, n_0_1595, n_0_1594, n_0_1593, n_0_1592, n_0_1591, 
      n_0_1590, n_0_1589, n_0_1588, n_0_1587, n_0_1586, n_0_1585, n_0_1584, 
      n_0_1583, n_0_1582, n_0_1581, n_0_1580, n_0_1579, n_0_1578, n_0_1577, 
      n_0_1576, n_0_1575, n_0_1574, n_0_1573, n_0_1572, n_0_1571, n_0_1570, 
      n_0_1569, n_0_1568}), .p_1({n_0_1662, n_0_1661, n_0_1660, n_0_1659, 
      n_0_1658, n_0_1657, n_0_1656, n_0_1655, n_0_1654, n_0_1653, n_0_1652, 
      n_0_1651, n_0_1650, n_0_1649, n_0_1648, n_0_1647, n_0_1646, n_0_1645, 
      n_0_1644, n_0_1643, n_0_1642, n_0_1641, n_0_1640, n_0_1639, n_0_1638, 
      n_0_1637, n_0_1636, n_0_1635, n_0_1634, n_0_1633, n_0_1632, n_0_1631}));
   INV_X1 i_0_68_0 (.A(multiplier2[17]), .ZN(n_0_68_0));
   AND2_X1 i_0_68_1 (.A1(n_0_68_0), .A2(multiplier2[16]), .ZN(n_0_1664));
   NOR2_X1 i_0_68_2 (.A1(n_0_68_0), .A2(multiplier2[16]), .ZN(n_0_1665));
   NOR2_X1 i_0_68_3 (.A1(n_0_1664), .A2(n_0_1665), .ZN(n_0_1663));
   AOI222_X1 i_0_69_0 (.A1(n_0_1631), .A2(n_0_1664), .B1(n_0_1599), .B2(n_0_1665), 
      .C1(n_0_1568), .C2(n_0_1663), .ZN(n_0_69_0));
   INV_X1 i_0_69_1 (.A(n_0_69_0), .ZN(product[17]));
   AOI222_X1 i_0_69_2 (.A1(n_0_1664), .A2(n_0_1632), .B1(n_0_1665), .B2(n_0_1600), 
      .C1(n_0_1663), .C2(n_0_1569), .ZN(n_0_69_1));
   INV_X1 i_0_69_3 (.A(n_0_69_1), .ZN(n_0_1666));
   AOI222_X1 i_0_69_4 (.A1(n_0_1664), .A2(n_0_1633), .B1(n_0_1665), .B2(n_0_1601), 
      .C1(n_0_1663), .C2(n_0_1570), .ZN(n_0_69_2));
   INV_X1 i_0_69_5 (.A(n_0_69_2), .ZN(n_0_1667));
   AOI222_X1 i_0_69_6 (.A1(n_0_1664), .A2(n_0_1634), .B1(n_0_1665), .B2(n_0_1602), 
      .C1(n_0_1663), .C2(n_0_1571), .ZN(n_0_69_3));
   INV_X1 i_0_69_7 (.A(n_0_69_3), .ZN(n_0_1668));
   AOI222_X1 i_0_69_8 (.A1(n_0_1664), .A2(n_0_1635), .B1(n_0_1665), .B2(n_0_1603), 
      .C1(n_0_1663), .C2(n_0_1572), .ZN(n_0_69_4));
   INV_X1 i_0_69_9 (.A(n_0_69_4), .ZN(n_0_1669));
   AOI222_X1 i_0_69_10 (.A1(n_0_1664), .A2(n_0_1636), .B1(n_0_1665), .B2(
      n_0_1604), .C1(n_0_1663), .C2(n_0_1573), .ZN(n_0_69_5));
   INV_X1 i_0_69_11 (.A(n_0_69_5), .ZN(n_0_1670));
   AOI222_X1 i_0_69_12 (.A1(n_0_1664), .A2(n_0_1637), .B1(n_0_1665), .B2(
      n_0_1605), .C1(n_0_1663), .C2(n_0_1574), .ZN(n_0_69_6));
   INV_X1 i_0_69_13 (.A(n_0_69_6), .ZN(n_0_1671));
   AOI222_X1 i_0_69_14 (.A1(n_0_1664), .A2(n_0_1638), .B1(n_0_1665), .B2(
      n_0_1606), .C1(n_0_1663), .C2(n_0_1575), .ZN(n_0_69_7));
   INV_X1 i_0_69_15 (.A(n_0_69_7), .ZN(n_0_1672));
   AOI222_X1 i_0_69_16 (.A1(n_0_1664), .A2(n_0_1639), .B1(n_0_1665), .B2(
      n_0_1607), .C1(n_0_1663), .C2(n_0_1576), .ZN(n_0_69_8));
   INV_X1 i_0_69_17 (.A(n_0_69_8), .ZN(n_0_1673));
   AOI222_X1 i_0_69_18 (.A1(n_0_1664), .A2(n_0_1640), .B1(n_0_1665), .B2(
      n_0_1608), .C1(n_0_1663), .C2(n_0_1577), .ZN(n_0_69_9));
   INV_X1 i_0_69_19 (.A(n_0_69_9), .ZN(n_0_1674));
   AOI222_X1 i_0_69_20 (.A1(n_0_1664), .A2(n_0_1641), .B1(n_0_1665), .B2(
      n_0_1609), .C1(n_0_1663), .C2(n_0_1578), .ZN(n_0_69_10));
   INV_X1 i_0_69_21 (.A(n_0_69_10), .ZN(n_0_1675));
   AOI222_X1 i_0_69_22 (.A1(n_0_1664), .A2(n_0_1642), .B1(n_0_1665), .B2(
      n_0_1610), .C1(n_0_1663), .C2(n_0_1579), .ZN(n_0_69_11));
   INV_X1 i_0_69_23 (.A(n_0_69_11), .ZN(n_0_1676));
   AOI222_X1 i_0_69_24 (.A1(n_0_1664), .A2(n_0_1643), .B1(n_0_1665), .B2(
      n_0_1611), .C1(n_0_1663), .C2(n_0_1580), .ZN(n_0_69_12));
   INV_X1 i_0_69_25 (.A(n_0_69_12), .ZN(n_0_1677));
   AOI222_X1 i_0_69_26 (.A1(n_0_1664), .A2(n_0_1644), .B1(n_0_1665), .B2(
      n_0_1612), .C1(n_0_1663), .C2(n_0_1581), .ZN(n_0_69_13));
   INV_X1 i_0_69_27 (.A(n_0_69_13), .ZN(n_0_1678));
   AOI222_X1 i_0_69_28 (.A1(n_0_1664), .A2(n_0_1645), .B1(n_0_1665), .B2(
      n_0_1613), .C1(n_0_1663), .C2(n_0_1582), .ZN(n_0_69_14));
   INV_X1 i_0_69_29 (.A(n_0_69_14), .ZN(n_0_1679));
   AOI222_X1 i_0_69_30 (.A1(n_0_1664), .A2(n_0_1646), .B1(n_0_1665), .B2(
      n_0_1614), .C1(n_0_1663), .C2(n_0_1583), .ZN(n_0_69_15));
   INV_X1 i_0_69_31 (.A(n_0_69_15), .ZN(n_0_1680));
   AOI222_X1 i_0_69_32 (.A1(n_0_1664), .A2(n_0_1647), .B1(n_0_1665), .B2(
      n_0_1615), .C1(n_0_1663), .C2(n_0_1584), .ZN(n_0_69_16));
   INV_X1 i_0_69_33 (.A(n_0_69_16), .ZN(n_0_1681));
   AOI222_X1 i_0_69_34 (.A1(n_0_1664), .A2(n_0_1648), .B1(n_0_1665), .B2(
      n_0_1616), .C1(n_0_1663), .C2(n_0_1585), .ZN(n_0_69_17));
   INV_X1 i_0_69_35 (.A(n_0_69_17), .ZN(n_0_1682));
   AOI222_X1 i_0_69_36 (.A1(n_0_1664), .A2(n_0_1649), .B1(n_0_1665), .B2(
      n_0_1617), .C1(n_0_1663), .C2(n_0_1586), .ZN(n_0_69_18));
   INV_X1 i_0_69_37 (.A(n_0_69_18), .ZN(n_0_1683));
   AOI222_X1 i_0_69_38 (.A1(n_0_1664), .A2(n_0_1650), .B1(n_0_1665), .B2(
      n_0_1618), .C1(n_0_1663), .C2(n_0_1587), .ZN(n_0_69_19));
   INV_X1 i_0_69_39 (.A(n_0_69_19), .ZN(n_0_1684));
   AOI222_X1 i_0_69_40 (.A1(n_0_1664), .A2(n_0_1651), .B1(n_0_1665), .B2(
      n_0_1619), .C1(n_0_1663), .C2(n_0_1588), .ZN(n_0_69_20));
   INV_X1 i_0_69_41 (.A(n_0_69_20), .ZN(n_0_1685));
   AOI222_X1 i_0_69_42 (.A1(n_0_1664), .A2(n_0_1652), .B1(n_0_1665), .B2(
      n_0_1620), .C1(n_0_1663), .C2(n_0_1589), .ZN(n_0_69_21));
   INV_X1 i_0_69_43 (.A(n_0_69_21), .ZN(n_0_1686));
   AOI222_X1 i_0_69_44 (.A1(n_0_1664), .A2(n_0_1653), .B1(n_0_1665), .B2(
      n_0_1621), .C1(n_0_1663), .C2(n_0_1590), .ZN(n_0_69_22));
   INV_X1 i_0_69_45 (.A(n_0_69_22), .ZN(n_0_1687));
   AOI222_X1 i_0_69_46 (.A1(n_0_1664), .A2(n_0_1654), .B1(n_0_1665), .B2(
      n_0_1622), .C1(n_0_1663), .C2(n_0_1591), .ZN(n_0_69_23));
   INV_X1 i_0_69_47 (.A(n_0_69_23), .ZN(n_0_1688));
   AOI222_X1 i_0_69_48 (.A1(n_0_1664), .A2(n_0_1655), .B1(n_0_1665), .B2(
      n_0_1623), .C1(n_0_1663), .C2(n_0_1592), .ZN(n_0_69_24));
   INV_X1 i_0_69_49 (.A(n_0_69_24), .ZN(n_0_1689));
   AOI222_X1 i_0_69_50 (.A1(n_0_1664), .A2(n_0_1656), .B1(n_0_1665), .B2(
      n_0_1624), .C1(n_0_1663), .C2(n_0_1593), .ZN(n_0_69_25));
   INV_X1 i_0_69_51 (.A(n_0_69_25), .ZN(n_0_1690));
   AOI222_X1 i_0_69_52 (.A1(n_0_1664), .A2(n_0_1657), .B1(n_0_1665), .B2(
      n_0_1625), .C1(n_0_1663), .C2(n_0_1594), .ZN(n_0_69_26));
   INV_X1 i_0_69_53 (.A(n_0_69_26), .ZN(n_0_1691));
   AOI222_X1 i_0_69_54 (.A1(n_0_1664), .A2(n_0_1658), .B1(n_0_1665), .B2(
      n_0_1626), .C1(n_0_1663), .C2(n_0_1595), .ZN(n_0_69_27));
   INV_X1 i_0_69_55 (.A(n_0_69_27), .ZN(n_0_1692));
   AOI222_X1 i_0_69_56 (.A1(n_0_1664), .A2(n_0_1659), .B1(n_0_1665), .B2(
      n_0_1627), .C1(n_0_1663), .C2(n_0_1596), .ZN(n_0_69_28));
   INV_X1 i_0_69_57 (.A(n_0_69_28), .ZN(n_0_1693));
   AOI222_X1 i_0_69_58 (.A1(n_0_1664), .A2(n_0_1660), .B1(n_0_1665), .B2(
      n_0_1628), .C1(n_0_1663), .C2(n_0_1597), .ZN(n_0_69_29));
   INV_X1 i_0_69_59 (.A(n_0_69_29), .ZN(n_0_1694));
   AND2_X1 i_0_69_60 (.A1(n_0_1663), .A2(n_0_1598), .ZN(n_0_69_30));
   AOI221_X1 i_0_69_61 (.A(n_0_69_30), .B1(n_0_1664), .B2(n_0_1661), .C1(
      n_0_1665), .C2(n_0_1629), .ZN(n_0_69_31));
   INV_X1 i_0_69_62 (.A(n_0_69_31), .ZN(n_0_1695));
   AOI221_X1 i_0_69_63 (.A(n_0_69_30), .B1(n_0_1664), .B2(n_0_1662), .C1(
      n_0_1665), .C2(n_0_1630), .ZN(n_0_69_32));
   INV_X1 i_0_69_64 (.A(n_0_69_32), .ZN(n_0_1696));
   datapath__0_68 i_0_70 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_35, 
      n_0_1696, n_0_1695, n_0_1694, n_0_1693, n_0_1692, n_0_1691, n_0_1690, 
      n_0_1689, n_0_1688, n_0_1687, n_0_1686, n_0_1685, n_0_1684, n_0_1683, 
      n_0_1682, n_0_1681, n_0_1680, n_0_1679, n_0_1678, n_0_1677, n_0_1676, 
      n_0_1675, n_0_1674, n_0_1673, n_0_1672, n_0_1671, n_0_1670, n_0_1669, 
      n_0_1668, n_0_1667, n_0_1666}), .p_2({n_0_1728, n_0_1727, n_0_1726, 
      n_0_1725, n_0_1724, n_0_1723, n_0_1722, n_0_1721, n_0_1720, n_0_1719, 
      n_0_1718, n_0_1717, n_0_1716, n_0_1715, n_0_1714, n_0_1713, n_0_1712, 
      n_0_1711, n_0_1710, n_0_1709, n_0_1708, n_0_1707, n_0_1706, n_0_1705, 
      n_0_1704, n_0_1703, n_0_1702, n_0_1701, n_0_1700, n_0_1699, n_0_1698, 
      n_0_1697}));
   datapath__0_69 i_0_71 (.multiplicand2(multiplicand2), .p_0({uc_36, n_0_1696, 
      n_0_1695, n_0_1694, n_0_1693, n_0_1692, n_0_1691, n_0_1690, n_0_1689, 
      n_0_1688, n_0_1687, n_0_1686, n_0_1685, n_0_1684, n_0_1683, n_0_1682, 
      n_0_1681, n_0_1680, n_0_1679, n_0_1678, n_0_1677, n_0_1676, n_0_1675, 
      n_0_1674, n_0_1673, n_0_1672, n_0_1671, n_0_1670, n_0_1669, n_0_1668, 
      n_0_1667, n_0_1666}), .p_1({n_0_1760, n_0_1759, n_0_1758, n_0_1757, 
      n_0_1756, n_0_1755, n_0_1754, n_0_1753, n_0_1752, n_0_1751, n_0_1750, 
      n_0_1749, n_0_1748, n_0_1747, n_0_1746, n_0_1745, n_0_1744, n_0_1743, 
      n_0_1742, n_0_1741, n_0_1740, n_0_1739, n_0_1738, n_0_1737, n_0_1736, 
      n_0_1735, n_0_1734, n_0_1733, n_0_1732, n_0_1731, n_0_1730, n_0_1729}));
   INV_X1 i_0_72_0 (.A(multiplier2[18]), .ZN(n_0_72_0));
   AND2_X1 i_0_72_1 (.A1(n_0_72_0), .A2(multiplier2[17]), .ZN(n_0_1762));
   NOR2_X1 i_0_72_2 (.A1(n_0_72_0), .A2(multiplier2[17]), .ZN(n_0_1763));
   NOR2_X1 i_0_72_3 (.A1(n_0_1762), .A2(n_0_1763), .ZN(n_0_1761));
   AOI222_X1 i_0_73_0 (.A1(n_0_1729), .A2(n_0_1762), .B1(n_0_1697), .B2(n_0_1763), 
      .C1(n_0_1666), .C2(n_0_1761), .ZN(n_0_73_0));
   INV_X1 i_0_73_1 (.A(n_0_73_0), .ZN(product[18]));
   AOI222_X1 i_0_73_2 (.A1(n_0_1762), .A2(n_0_1730), .B1(n_0_1763), .B2(n_0_1698), 
      .C1(n_0_1761), .C2(n_0_1667), .ZN(n_0_73_1));
   INV_X1 i_0_73_3 (.A(n_0_73_1), .ZN(n_0_1764));
   AOI222_X1 i_0_73_4 (.A1(n_0_1762), .A2(n_0_1731), .B1(n_0_1763), .B2(n_0_1699), 
      .C1(n_0_1761), .C2(n_0_1668), .ZN(n_0_73_2));
   INV_X1 i_0_73_5 (.A(n_0_73_2), .ZN(n_0_1765));
   AOI222_X1 i_0_73_6 (.A1(n_0_1762), .A2(n_0_1732), .B1(n_0_1763), .B2(n_0_1700), 
      .C1(n_0_1761), .C2(n_0_1669), .ZN(n_0_73_3));
   INV_X1 i_0_73_7 (.A(n_0_73_3), .ZN(n_0_1766));
   AOI222_X1 i_0_73_8 (.A1(n_0_1762), .A2(n_0_1733), .B1(n_0_1763), .B2(n_0_1701), 
      .C1(n_0_1761), .C2(n_0_1670), .ZN(n_0_73_4));
   INV_X1 i_0_73_9 (.A(n_0_73_4), .ZN(n_0_1767));
   AOI222_X1 i_0_73_10 (.A1(n_0_1762), .A2(n_0_1734), .B1(n_0_1763), .B2(
      n_0_1702), .C1(n_0_1761), .C2(n_0_1671), .ZN(n_0_73_5));
   INV_X1 i_0_73_11 (.A(n_0_73_5), .ZN(n_0_1768));
   AOI222_X1 i_0_73_12 (.A1(n_0_1762), .A2(n_0_1735), .B1(n_0_1763), .B2(
      n_0_1703), .C1(n_0_1761), .C2(n_0_1672), .ZN(n_0_73_6));
   INV_X1 i_0_73_13 (.A(n_0_73_6), .ZN(n_0_1769));
   AOI222_X1 i_0_73_14 (.A1(n_0_1762), .A2(n_0_1736), .B1(n_0_1763), .B2(
      n_0_1704), .C1(n_0_1761), .C2(n_0_1673), .ZN(n_0_73_7));
   INV_X1 i_0_73_15 (.A(n_0_73_7), .ZN(n_0_1770));
   AOI222_X1 i_0_73_16 (.A1(n_0_1762), .A2(n_0_1737), .B1(n_0_1763), .B2(
      n_0_1705), .C1(n_0_1761), .C2(n_0_1674), .ZN(n_0_73_8));
   INV_X1 i_0_73_17 (.A(n_0_73_8), .ZN(n_0_1771));
   AOI222_X1 i_0_73_18 (.A1(n_0_1762), .A2(n_0_1738), .B1(n_0_1763), .B2(
      n_0_1706), .C1(n_0_1761), .C2(n_0_1675), .ZN(n_0_73_9));
   INV_X1 i_0_73_19 (.A(n_0_73_9), .ZN(n_0_1772));
   AOI222_X1 i_0_73_20 (.A1(n_0_1762), .A2(n_0_1739), .B1(n_0_1763), .B2(
      n_0_1707), .C1(n_0_1761), .C2(n_0_1676), .ZN(n_0_73_10));
   INV_X1 i_0_73_21 (.A(n_0_73_10), .ZN(n_0_1773));
   AOI222_X1 i_0_73_22 (.A1(n_0_1762), .A2(n_0_1740), .B1(n_0_1763), .B2(
      n_0_1708), .C1(n_0_1761), .C2(n_0_1677), .ZN(n_0_73_11));
   INV_X1 i_0_73_23 (.A(n_0_73_11), .ZN(n_0_1774));
   AOI222_X1 i_0_73_24 (.A1(n_0_1762), .A2(n_0_1741), .B1(n_0_1763), .B2(
      n_0_1709), .C1(n_0_1761), .C2(n_0_1678), .ZN(n_0_73_12));
   INV_X1 i_0_73_25 (.A(n_0_73_12), .ZN(n_0_1775));
   AOI222_X1 i_0_73_26 (.A1(n_0_1762), .A2(n_0_1742), .B1(n_0_1763), .B2(
      n_0_1710), .C1(n_0_1761), .C2(n_0_1679), .ZN(n_0_73_13));
   INV_X1 i_0_73_27 (.A(n_0_73_13), .ZN(n_0_1776));
   AOI222_X1 i_0_73_28 (.A1(n_0_1762), .A2(n_0_1743), .B1(n_0_1763), .B2(
      n_0_1711), .C1(n_0_1761), .C2(n_0_1680), .ZN(n_0_73_14));
   INV_X1 i_0_73_29 (.A(n_0_73_14), .ZN(n_0_1777));
   AOI222_X1 i_0_73_30 (.A1(n_0_1762), .A2(n_0_1744), .B1(n_0_1763), .B2(
      n_0_1712), .C1(n_0_1761), .C2(n_0_1681), .ZN(n_0_73_15));
   INV_X1 i_0_73_31 (.A(n_0_73_15), .ZN(n_0_1778));
   AOI222_X1 i_0_73_32 (.A1(n_0_1762), .A2(n_0_1745), .B1(n_0_1763), .B2(
      n_0_1713), .C1(n_0_1761), .C2(n_0_1682), .ZN(n_0_73_16));
   INV_X1 i_0_73_33 (.A(n_0_73_16), .ZN(n_0_1779));
   AOI222_X1 i_0_73_34 (.A1(n_0_1762), .A2(n_0_1746), .B1(n_0_1763), .B2(
      n_0_1714), .C1(n_0_1761), .C2(n_0_1683), .ZN(n_0_73_17));
   INV_X1 i_0_73_35 (.A(n_0_73_17), .ZN(n_0_1780));
   AOI222_X1 i_0_73_36 (.A1(n_0_1762), .A2(n_0_1747), .B1(n_0_1763), .B2(
      n_0_1715), .C1(n_0_1761), .C2(n_0_1684), .ZN(n_0_73_18));
   INV_X1 i_0_73_37 (.A(n_0_73_18), .ZN(n_0_1781));
   AOI222_X1 i_0_73_38 (.A1(n_0_1762), .A2(n_0_1748), .B1(n_0_1763), .B2(
      n_0_1716), .C1(n_0_1761), .C2(n_0_1685), .ZN(n_0_73_19));
   INV_X1 i_0_73_39 (.A(n_0_73_19), .ZN(n_0_1782));
   AOI222_X1 i_0_73_40 (.A1(n_0_1762), .A2(n_0_1749), .B1(n_0_1763), .B2(
      n_0_1717), .C1(n_0_1761), .C2(n_0_1686), .ZN(n_0_73_20));
   INV_X1 i_0_73_41 (.A(n_0_73_20), .ZN(n_0_1783));
   AOI222_X1 i_0_73_42 (.A1(n_0_1762), .A2(n_0_1750), .B1(n_0_1763), .B2(
      n_0_1718), .C1(n_0_1761), .C2(n_0_1687), .ZN(n_0_73_21));
   INV_X1 i_0_73_43 (.A(n_0_73_21), .ZN(n_0_1784));
   AOI222_X1 i_0_73_44 (.A1(n_0_1762), .A2(n_0_1751), .B1(n_0_1763), .B2(
      n_0_1719), .C1(n_0_1761), .C2(n_0_1688), .ZN(n_0_73_22));
   INV_X1 i_0_73_45 (.A(n_0_73_22), .ZN(n_0_1785));
   AOI222_X1 i_0_73_46 (.A1(n_0_1762), .A2(n_0_1752), .B1(n_0_1763), .B2(
      n_0_1720), .C1(n_0_1761), .C2(n_0_1689), .ZN(n_0_73_23));
   INV_X1 i_0_73_47 (.A(n_0_73_23), .ZN(n_0_1786));
   AOI222_X1 i_0_73_48 (.A1(n_0_1762), .A2(n_0_1753), .B1(n_0_1763), .B2(
      n_0_1721), .C1(n_0_1761), .C2(n_0_1690), .ZN(n_0_73_24));
   INV_X1 i_0_73_49 (.A(n_0_73_24), .ZN(n_0_1787));
   AOI222_X1 i_0_73_50 (.A1(n_0_1762), .A2(n_0_1754), .B1(n_0_1763), .B2(
      n_0_1722), .C1(n_0_1761), .C2(n_0_1691), .ZN(n_0_73_25));
   INV_X1 i_0_73_51 (.A(n_0_73_25), .ZN(n_0_1788));
   AOI222_X1 i_0_73_52 (.A1(n_0_1762), .A2(n_0_1755), .B1(n_0_1763), .B2(
      n_0_1723), .C1(n_0_1761), .C2(n_0_1692), .ZN(n_0_73_26));
   INV_X1 i_0_73_53 (.A(n_0_73_26), .ZN(n_0_1789));
   AOI222_X1 i_0_73_54 (.A1(n_0_1762), .A2(n_0_1756), .B1(n_0_1763), .B2(
      n_0_1724), .C1(n_0_1761), .C2(n_0_1693), .ZN(n_0_73_27));
   INV_X1 i_0_73_55 (.A(n_0_73_27), .ZN(n_0_1790));
   AOI222_X1 i_0_73_56 (.A1(n_0_1762), .A2(n_0_1757), .B1(n_0_1763), .B2(
      n_0_1725), .C1(n_0_1761), .C2(n_0_1694), .ZN(n_0_73_28));
   INV_X1 i_0_73_57 (.A(n_0_73_28), .ZN(n_0_1791));
   AOI222_X1 i_0_73_58 (.A1(n_0_1762), .A2(n_0_1758), .B1(n_0_1763), .B2(
      n_0_1726), .C1(n_0_1761), .C2(n_0_1695), .ZN(n_0_73_29));
   INV_X1 i_0_73_59 (.A(n_0_73_29), .ZN(n_0_1792));
   AND2_X1 i_0_73_60 (.A1(n_0_1761), .A2(n_0_1696), .ZN(n_0_73_30));
   AOI221_X1 i_0_73_61 (.A(n_0_73_30), .B1(n_0_1762), .B2(n_0_1759), .C1(
      n_0_1763), .C2(n_0_1727), .ZN(n_0_73_31));
   INV_X1 i_0_73_62 (.A(n_0_73_31), .ZN(n_0_1793));
   AOI221_X1 i_0_73_63 (.A(n_0_73_30), .B1(n_0_1762), .B2(n_0_1760), .C1(
      n_0_1763), .C2(n_0_1728), .ZN(n_0_73_32));
   INV_X1 i_0_73_64 (.A(n_0_73_32), .ZN(n_0_1794));
   datapath__0_72 i_0_74 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_37, 
      n_0_1794, n_0_1793, n_0_1792, n_0_1791, n_0_1790, n_0_1789, n_0_1788, 
      n_0_1787, n_0_1786, n_0_1785, n_0_1784, n_0_1783, n_0_1782, n_0_1781, 
      n_0_1780, n_0_1779, n_0_1778, n_0_1777, n_0_1776, n_0_1775, n_0_1774, 
      n_0_1773, n_0_1772, n_0_1771, n_0_1770, n_0_1769, n_0_1768, n_0_1767, 
      n_0_1766, n_0_1765, n_0_1764}), .p_2({n_0_1826, n_0_1825, n_0_1824, 
      n_0_1823, n_0_1822, n_0_1821, n_0_1820, n_0_1819, n_0_1818, n_0_1817, 
      n_0_1816, n_0_1815, n_0_1814, n_0_1813, n_0_1812, n_0_1811, n_0_1810, 
      n_0_1809, n_0_1808, n_0_1807, n_0_1806, n_0_1805, n_0_1804, n_0_1803, 
      n_0_1802, n_0_1801, n_0_1800, n_0_1799, n_0_1798, n_0_1797, n_0_1796, 
      n_0_1795}));
   datapath__0_73 i_0_75 (.multiplicand2(multiplicand2), .p_0({uc_38, n_0_1794, 
      n_0_1793, n_0_1792, n_0_1791, n_0_1790, n_0_1789, n_0_1788, n_0_1787, 
      n_0_1786, n_0_1785, n_0_1784, n_0_1783, n_0_1782, n_0_1781, n_0_1780, 
      n_0_1779, n_0_1778, n_0_1777, n_0_1776, n_0_1775, n_0_1774, n_0_1773, 
      n_0_1772, n_0_1771, n_0_1770, n_0_1769, n_0_1768, n_0_1767, n_0_1766, 
      n_0_1765, n_0_1764}), .p_1({n_0_1858, n_0_1857, n_0_1856, n_0_1855, 
      n_0_1854, n_0_1853, n_0_1852, n_0_1851, n_0_1850, n_0_1849, n_0_1848, 
      n_0_1847, n_0_1846, n_0_1845, n_0_1844, n_0_1843, n_0_1842, n_0_1841, 
      n_0_1840, n_0_1839, n_0_1838, n_0_1837, n_0_1836, n_0_1835, n_0_1834, 
      n_0_1833, n_0_1832, n_0_1831, n_0_1830, n_0_1829, n_0_1828, n_0_1827}));
   INV_X1 i_0_76_0 (.A(multiplier2[19]), .ZN(n_0_76_0));
   AND2_X1 i_0_76_1 (.A1(n_0_76_0), .A2(multiplier2[18]), .ZN(n_0_1860));
   NOR2_X1 i_0_76_2 (.A1(n_0_76_0), .A2(multiplier2[18]), .ZN(n_0_1861));
   NOR2_X1 i_0_76_3 (.A1(n_0_1860), .A2(n_0_1861), .ZN(n_0_1859));
   AOI222_X1 i_0_77_0 (.A1(n_0_1827), .A2(n_0_1860), .B1(n_0_1795), .B2(n_0_1861), 
      .C1(n_0_1764), .C2(n_0_1859), .ZN(n_0_77_0));
   INV_X1 i_0_77_1 (.A(n_0_77_0), .ZN(product[19]));
   AOI222_X1 i_0_77_2 (.A1(n_0_1860), .A2(n_0_1828), .B1(n_0_1861), .B2(n_0_1796), 
      .C1(n_0_1859), .C2(n_0_1765), .ZN(n_0_77_1));
   INV_X1 i_0_77_3 (.A(n_0_77_1), .ZN(n_0_1862));
   AOI222_X1 i_0_77_4 (.A1(n_0_1860), .A2(n_0_1829), .B1(n_0_1861), .B2(n_0_1797), 
      .C1(n_0_1859), .C2(n_0_1766), .ZN(n_0_77_2));
   INV_X1 i_0_77_5 (.A(n_0_77_2), .ZN(n_0_1863));
   AOI222_X1 i_0_77_6 (.A1(n_0_1860), .A2(n_0_1830), .B1(n_0_1861), .B2(n_0_1798), 
      .C1(n_0_1859), .C2(n_0_1767), .ZN(n_0_77_3));
   INV_X1 i_0_77_7 (.A(n_0_77_3), .ZN(n_0_1864));
   AOI222_X1 i_0_77_8 (.A1(n_0_1860), .A2(n_0_1831), .B1(n_0_1861), .B2(n_0_1799), 
      .C1(n_0_1859), .C2(n_0_1768), .ZN(n_0_77_4));
   INV_X1 i_0_77_9 (.A(n_0_77_4), .ZN(n_0_1865));
   AOI222_X1 i_0_77_10 (.A1(n_0_1860), .A2(n_0_1832), .B1(n_0_1861), .B2(
      n_0_1800), .C1(n_0_1859), .C2(n_0_1769), .ZN(n_0_77_5));
   INV_X1 i_0_77_11 (.A(n_0_77_5), .ZN(n_0_1866));
   AOI222_X1 i_0_77_12 (.A1(n_0_1860), .A2(n_0_1833), .B1(n_0_1861), .B2(
      n_0_1801), .C1(n_0_1859), .C2(n_0_1770), .ZN(n_0_77_6));
   INV_X1 i_0_77_13 (.A(n_0_77_6), .ZN(n_0_1867));
   AOI222_X1 i_0_77_14 (.A1(n_0_1860), .A2(n_0_1834), .B1(n_0_1861), .B2(
      n_0_1802), .C1(n_0_1859), .C2(n_0_1771), .ZN(n_0_77_7));
   INV_X1 i_0_77_15 (.A(n_0_77_7), .ZN(n_0_1868));
   AOI222_X1 i_0_77_16 (.A1(n_0_1860), .A2(n_0_1835), .B1(n_0_1861), .B2(
      n_0_1803), .C1(n_0_1859), .C2(n_0_1772), .ZN(n_0_77_8));
   INV_X1 i_0_77_17 (.A(n_0_77_8), .ZN(n_0_1869));
   AOI222_X1 i_0_77_18 (.A1(n_0_1860), .A2(n_0_1836), .B1(n_0_1861), .B2(
      n_0_1804), .C1(n_0_1859), .C2(n_0_1773), .ZN(n_0_77_9));
   INV_X1 i_0_77_19 (.A(n_0_77_9), .ZN(n_0_1870));
   AOI222_X1 i_0_77_20 (.A1(n_0_1860), .A2(n_0_1837), .B1(n_0_1861), .B2(
      n_0_1805), .C1(n_0_1859), .C2(n_0_1774), .ZN(n_0_77_10));
   INV_X1 i_0_77_21 (.A(n_0_77_10), .ZN(n_0_1871));
   AOI222_X1 i_0_77_22 (.A1(n_0_1860), .A2(n_0_1838), .B1(n_0_1861), .B2(
      n_0_1806), .C1(n_0_1859), .C2(n_0_1775), .ZN(n_0_77_11));
   INV_X1 i_0_77_23 (.A(n_0_77_11), .ZN(n_0_1872));
   AOI222_X1 i_0_77_24 (.A1(n_0_1860), .A2(n_0_1839), .B1(n_0_1861), .B2(
      n_0_1807), .C1(n_0_1859), .C2(n_0_1776), .ZN(n_0_77_12));
   INV_X1 i_0_77_25 (.A(n_0_77_12), .ZN(n_0_1873));
   AOI222_X1 i_0_77_26 (.A1(n_0_1860), .A2(n_0_1840), .B1(n_0_1861), .B2(
      n_0_1808), .C1(n_0_1859), .C2(n_0_1777), .ZN(n_0_77_13));
   INV_X1 i_0_77_27 (.A(n_0_77_13), .ZN(n_0_1874));
   AOI222_X1 i_0_77_28 (.A1(n_0_1860), .A2(n_0_1841), .B1(n_0_1861), .B2(
      n_0_1809), .C1(n_0_1859), .C2(n_0_1778), .ZN(n_0_77_14));
   INV_X1 i_0_77_29 (.A(n_0_77_14), .ZN(n_0_1875));
   AOI222_X1 i_0_77_30 (.A1(n_0_1860), .A2(n_0_1842), .B1(n_0_1861), .B2(
      n_0_1810), .C1(n_0_1859), .C2(n_0_1779), .ZN(n_0_77_15));
   INV_X1 i_0_77_31 (.A(n_0_77_15), .ZN(n_0_1876));
   AOI222_X1 i_0_77_32 (.A1(n_0_1860), .A2(n_0_1843), .B1(n_0_1861), .B2(
      n_0_1811), .C1(n_0_1859), .C2(n_0_1780), .ZN(n_0_77_16));
   INV_X1 i_0_77_33 (.A(n_0_77_16), .ZN(n_0_1877));
   AOI222_X1 i_0_77_34 (.A1(n_0_1860), .A2(n_0_1844), .B1(n_0_1861), .B2(
      n_0_1812), .C1(n_0_1859), .C2(n_0_1781), .ZN(n_0_77_17));
   INV_X1 i_0_77_35 (.A(n_0_77_17), .ZN(n_0_1878));
   AOI222_X1 i_0_77_36 (.A1(n_0_1860), .A2(n_0_1845), .B1(n_0_1861), .B2(
      n_0_1813), .C1(n_0_1859), .C2(n_0_1782), .ZN(n_0_77_18));
   INV_X1 i_0_77_37 (.A(n_0_77_18), .ZN(n_0_1879));
   AOI222_X1 i_0_77_38 (.A1(n_0_1860), .A2(n_0_1846), .B1(n_0_1861), .B2(
      n_0_1814), .C1(n_0_1859), .C2(n_0_1783), .ZN(n_0_77_19));
   INV_X1 i_0_77_39 (.A(n_0_77_19), .ZN(n_0_1880));
   AOI222_X1 i_0_77_40 (.A1(n_0_1860), .A2(n_0_1847), .B1(n_0_1861), .B2(
      n_0_1815), .C1(n_0_1859), .C2(n_0_1784), .ZN(n_0_77_20));
   INV_X1 i_0_77_41 (.A(n_0_77_20), .ZN(n_0_1881));
   AOI222_X1 i_0_77_42 (.A1(n_0_1860), .A2(n_0_1848), .B1(n_0_1861), .B2(
      n_0_1816), .C1(n_0_1859), .C2(n_0_1785), .ZN(n_0_77_21));
   INV_X1 i_0_77_43 (.A(n_0_77_21), .ZN(n_0_1882));
   AOI222_X1 i_0_77_44 (.A1(n_0_1860), .A2(n_0_1849), .B1(n_0_1861), .B2(
      n_0_1817), .C1(n_0_1859), .C2(n_0_1786), .ZN(n_0_77_22));
   INV_X1 i_0_77_45 (.A(n_0_77_22), .ZN(n_0_1883));
   AOI222_X1 i_0_77_46 (.A1(n_0_1860), .A2(n_0_1850), .B1(n_0_1861), .B2(
      n_0_1818), .C1(n_0_1859), .C2(n_0_1787), .ZN(n_0_77_23));
   INV_X1 i_0_77_47 (.A(n_0_77_23), .ZN(n_0_1884));
   AOI222_X1 i_0_77_48 (.A1(n_0_1860), .A2(n_0_1851), .B1(n_0_1861), .B2(
      n_0_1819), .C1(n_0_1859), .C2(n_0_1788), .ZN(n_0_77_24));
   INV_X1 i_0_77_49 (.A(n_0_77_24), .ZN(n_0_1885));
   AOI222_X1 i_0_77_50 (.A1(n_0_1860), .A2(n_0_1852), .B1(n_0_1861), .B2(
      n_0_1820), .C1(n_0_1859), .C2(n_0_1789), .ZN(n_0_77_25));
   INV_X1 i_0_77_51 (.A(n_0_77_25), .ZN(n_0_1886));
   AOI222_X1 i_0_77_52 (.A1(n_0_1860), .A2(n_0_1853), .B1(n_0_1861), .B2(
      n_0_1821), .C1(n_0_1859), .C2(n_0_1790), .ZN(n_0_77_26));
   INV_X1 i_0_77_53 (.A(n_0_77_26), .ZN(n_0_1887));
   AOI222_X1 i_0_77_54 (.A1(n_0_1860), .A2(n_0_1854), .B1(n_0_1861), .B2(
      n_0_1822), .C1(n_0_1859), .C2(n_0_1791), .ZN(n_0_77_27));
   INV_X1 i_0_77_55 (.A(n_0_77_27), .ZN(n_0_1888));
   AOI222_X1 i_0_77_56 (.A1(n_0_1860), .A2(n_0_1855), .B1(n_0_1861), .B2(
      n_0_1823), .C1(n_0_1859), .C2(n_0_1792), .ZN(n_0_77_28));
   INV_X1 i_0_77_57 (.A(n_0_77_28), .ZN(n_0_1889));
   AOI222_X1 i_0_77_58 (.A1(n_0_1860), .A2(n_0_1856), .B1(n_0_1861), .B2(
      n_0_1824), .C1(n_0_1859), .C2(n_0_1793), .ZN(n_0_77_29));
   INV_X1 i_0_77_59 (.A(n_0_77_29), .ZN(n_0_1890));
   AND2_X1 i_0_77_60 (.A1(n_0_1859), .A2(n_0_1794), .ZN(n_0_77_30));
   AOI221_X1 i_0_77_61 (.A(n_0_77_30), .B1(n_0_1860), .B2(n_0_1857), .C1(
      n_0_1861), .C2(n_0_1825), .ZN(n_0_77_31));
   INV_X1 i_0_77_62 (.A(n_0_77_31), .ZN(n_0_1891));
   AOI221_X1 i_0_77_63 (.A(n_0_77_30), .B1(n_0_1860), .B2(n_0_1858), .C1(
      n_0_1861), .C2(n_0_1826), .ZN(n_0_77_32));
   INV_X1 i_0_77_64 (.A(n_0_77_32), .ZN(n_0_1892));
   datapath__0_76 i_0_78 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_39, 
      n_0_1892, n_0_1891, n_0_1890, n_0_1889, n_0_1888, n_0_1887, n_0_1886, 
      n_0_1885, n_0_1884, n_0_1883, n_0_1882, n_0_1881, n_0_1880, n_0_1879, 
      n_0_1878, n_0_1877, n_0_1876, n_0_1875, n_0_1874, n_0_1873, n_0_1872, 
      n_0_1871, n_0_1870, n_0_1869, n_0_1868, n_0_1867, n_0_1866, n_0_1865, 
      n_0_1864, n_0_1863, n_0_1862}), .p_2({n_0_1924, n_0_1923, n_0_1922, 
      n_0_1921, n_0_1920, n_0_1919, n_0_1918, n_0_1917, n_0_1916, n_0_1915, 
      n_0_1914, n_0_1913, n_0_1912, n_0_1911, n_0_1910, n_0_1909, n_0_1908, 
      n_0_1907, n_0_1906, n_0_1905, n_0_1904, n_0_1903, n_0_1902, n_0_1901, 
      n_0_1900, n_0_1899, n_0_1898, n_0_1897, n_0_1896, n_0_1895, n_0_1894, 
      n_0_1893}));
   datapath__0_77 i_0_79 (.multiplicand2(multiplicand2), .p_0({uc_40, n_0_1892, 
      n_0_1891, n_0_1890, n_0_1889, n_0_1888, n_0_1887, n_0_1886, n_0_1885, 
      n_0_1884, n_0_1883, n_0_1882, n_0_1881, n_0_1880, n_0_1879, n_0_1878, 
      n_0_1877, n_0_1876, n_0_1875, n_0_1874, n_0_1873, n_0_1872, n_0_1871, 
      n_0_1870, n_0_1869, n_0_1868, n_0_1867, n_0_1866, n_0_1865, n_0_1864, 
      n_0_1863, n_0_1862}), .p_1({n_0_1956, n_0_1955, n_0_1954, n_0_1953, 
      n_0_1952, n_0_1951, n_0_1950, n_0_1949, n_0_1948, n_0_1947, n_0_1946, 
      n_0_1945, n_0_1944, n_0_1943, n_0_1942, n_0_1941, n_0_1940, n_0_1939, 
      n_0_1938, n_0_1937, n_0_1936, n_0_1935, n_0_1934, n_0_1933, n_0_1932, 
      n_0_1931, n_0_1930, n_0_1929, n_0_1928, n_0_1927, n_0_1926, n_0_1925}));
   INV_X1 i_0_80_0 (.A(multiplier2[20]), .ZN(n_0_80_0));
   AND2_X1 i_0_80_1 (.A1(n_0_80_0), .A2(multiplier2[19]), .ZN(n_0_1958));
   NOR2_X1 i_0_80_2 (.A1(n_0_80_0), .A2(multiplier2[19]), .ZN(n_0_1959));
   NOR2_X1 i_0_80_3 (.A1(n_0_1958), .A2(n_0_1959), .ZN(n_0_1957));
   AOI222_X1 i_0_81_0 (.A1(n_0_1925), .A2(n_0_1958), .B1(n_0_1893), .B2(n_0_1959), 
      .C1(n_0_1862), .C2(n_0_1957), .ZN(n_0_81_0));
   INV_X1 i_0_81_1 (.A(n_0_81_0), .ZN(product[20]));
   AOI222_X1 i_0_81_2 (.A1(n_0_1958), .A2(n_0_1926), .B1(n_0_1959), .B2(n_0_1894), 
      .C1(n_0_1957), .C2(n_0_1863), .ZN(n_0_81_1));
   INV_X1 i_0_81_3 (.A(n_0_81_1), .ZN(n_0_1960));
   AOI222_X1 i_0_81_4 (.A1(n_0_1958), .A2(n_0_1927), .B1(n_0_1959), .B2(n_0_1895), 
      .C1(n_0_1957), .C2(n_0_1864), .ZN(n_0_81_2));
   INV_X1 i_0_81_5 (.A(n_0_81_2), .ZN(n_0_1961));
   AOI222_X1 i_0_81_6 (.A1(n_0_1958), .A2(n_0_1928), .B1(n_0_1959), .B2(n_0_1896), 
      .C1(n_0_1957), .C2(n_0_1865), .ZN(n_0_81_3));
   INV_X1 i_0_81_7 (.A(n_0_81_3), .ZN(n_0_1962));
   AOI222_X1 i_0_81_8 (.A1(n_0_1958), .A2(n_0_1929), .B1(n_0_1959), .B2(n_0_1897), 
      .C1(n_0_1957), .C2(n_0_1866), .ZN(n_0_81_4));
   INV_X1 i_0_81_9 (.A(n_0_81_4), .ZN(n_0_1963));
   AOI222_X1 i_0_81_10 (.A1(n_0_1958), .A2(n_0_1930), .B1(n_0_1959), .B2(
      n_0_1898), .C1(n_0_1957), .C2(n_0_1867), .ZN(n_0_81_5));
   INV_X1 i_0_81_11 (.A(n_0_81_5), .ZN(n_0_1964));
   AOI222_X1 i_0_81_12 (.A1(n_0_1958), .A2(n_0_1931), .B1(n_0_1959), .B2(
      n_0_1899), .C1(n_0_1957), .C2(n_0_1868), .ZN(n_0_81_6));
   INV_X1 i_0_81_13 (.A(n_0_81_6), .ZN(n_0_1965));
   AOI222_X1 i_0_81_14 (.A1(n_0_1958), .A2(n_0_1932), .B1(n_0_1959), .B2(
      n_0_1900), .C1(n_0_1957), .C2(n_0_1869), .ZN(n_0_81_7));
   INV_X1 i_0_81_15 (.A(n_0_81_7), .ZN(n_0_1966));
   AOI222_X1 i_0_81_16 (.A1(n_0_1958), .A2(n_0_1933), .B1(n_0_1959), .B2(
      n_0_1901), .C1(n_0_1957), .C2(n_0_1870), .ZN(n_0_81_8));
   INV_X1 i_0_81_17 (.A(n_0_81_8), .ZN(n_0_1967));
   AOI222_X1 i_0_81_18 (.A1(n_0_1958), .A2(n_0_1934), .B1(n_0_1959), .B2(
      n_0_1902), .C1(n_0_1957), .C2(n_0_1871), .ZN(n_0_81_9));
   INV_X1 i_0_81_19 (.A(n_0_81_9), .ZN(n_0_1968));
   AOI222_X1 i_0_81_20 (.A1(n_0_1958), .A2(n_0_1935), .B1(n_0_1959), .B2(
      n_0_1903), .C1(n_0_1957), .C2(n_0_1872), .ZN(n_0_81_10));
   INV_X1 i_0_81_21 (.A(n_0_81_10), .ZN(n_0_1969));
   AOI222_X1 i_0_81_22 (.A1(n_0_1958), .A2(n_0_1936), .B1(n_0_1959), .B2(
      n_0_1904), .C1(n_0_1957), .C2(n_0_1873), .ZN(n_0_81_11));
   INV_X1 i_0_81_23 (.A(n_0_81_11), .ZN(n_0_1970));
   AOI222_X1 i_0_81_24 (.A1(n_0_1958), .A2(n_0_1937), .B1(n_0_1959), .B2(
      n_0_1905), .C1(n_0_1957), .C2(n_0_1874), .ZN(n_0_81_12));
   INV_X1 i_0_81_25 (.A(n_0_81_12), .ZN(n_0_1971));
   AOI222_X1 i_0_81_26 (.A1(n_0_1958), .A2(n_0_1938), .B1(n_0_1959), .B2(
      n_0_1906), .C1(n_0_1957), .C2(n_0_1875), .ZN(n_0_81_13));
   INV_X1 i_0_81_27 (.A(n_0_81_13), .ZN(n_0_1972));
   AOI222_X1 i_0_81_28 (.A1(n_0_1958), .A2(n_0_1939), .B1(n_0_1959), .B2(
      n_0_1907), .C1(n_0_1957), .C2(n_0_1876), .ZN(n_0_81_14));
   INV_X1 i_0_81_29 (.A(n_0_81_14), .ZN(n_0_1973));
   AOI222_X1 i_0_81_30 (.A1(n_0_1958), .A2(n_0_1940), .B1(n_0_1959), .B2(
      n_0_1908), .C1(n_0_1957), .C2(n_0_1877), .ZN(n_0_81_15));
   INV_X1 i_0_81_31 (.A(n_0_81_15), .ZN(n_0_1974));
   AOI222_X1 i_0_81_32 (.A1(n_0_1958), .A2(n_0_1941), .B1(n_0_1959), .B2(
      n_0_1909), .C1(n_0_1957), .C2(n_0_1878), .ZN(n_0_81_16));
   INV_X1 i_0_81_33 (.A(n_0_81_16), .ZN(n_0_1975));
   AOI222_X1 i_0_81_34 (.A1(n_0_1958), .A2(n_0_1942), .B1(n_0_1959), .B2(
      n_0_1910), .C1(n_0_1957), .C2(n_0_1879), .ZN(n_0_81_17));
   INV_X1 i_0_81_35 (.A(n_0_81_17), .ZN(n_0_1976));
   AOI222_X1 i_0_81_36 (.A1(n_0_1958), .A2(n_0_1943), .B1(n_0_1959), .B2(
      n_0_1911), .C1(n_0_1957), .C2(n_0_1880), .ZN(n_0_81_18));
   INV_X1 i_0_81_37 (.A(n_0_81_18), .ZN(n_0_1977));
   AOI222_X1 i_0_81_38 (.A1(n_0_1958), .A2(n_0_1944), .B1(n_0_1959), .B2(
      n_0_1912), .C1(n_0_1957), .C2(n_0_1881), .ZN(n_0_81_19));
   INV_X1 i_0_81_39 (.A(n_0_81_19), .ZN(n_0_1978));
   AOI222_X1 i_0_81_40 (.A1(n_0_1958), .A2(n_0_1945), .B1(n_0_1959), .B2(
      n_0_1913), .C1(n_0_1957), .C2(n_0_1882), .ZN(n_0_81_20));
   INV_X1 i_0_81_41 (.A(n_0_81_20), .ZN(n_0_1979));
   AOI222_X1 i_0_81_42 (.A1(n_0_1958), .A2(n_0_1946), .B1(n_0_1959), .B2(
      n_0_1914), .C1(n_0_1957), .C2(n_0_1883), .ZN(n_0_81_21));
   INV_X1 i_0_81_43 (.A(n_0_81_21), .ZN(n_0_1980));
   AOI222_X1 i_0_81_44 (.A1(n_0_1958), .A2(n_0_1947), .B1(n_0_1959), .B2(
      n_0_1915), .C1(n_0_1957), .C2(n_0_1884), .ZN(n_0_81_22));
   INV_X1 i_0_81_45 (.A(n_0_81_22), .ZN(n_0_1981));
   AOI222_X1 i_0_81_46 (.A1(n_0_1958), .A2(n_0_1948), .B1(n_0_1959), .B2(
      n_0_1916), .C1(n_0_1957), .C2(n_0_1885), .ZN(n_0_81_23));
   INV_X1 i_0_81_47 (.A(n_0_81_23), .ZN(n_0_1982));
   AOI222_X1 i_0_81_48 (.A1(n_0_1958), .A2(n_0_1949), .B1(n_0_1959), .B2(
      n_0_1917), .C1(n_0_1957), .C2(n_0_1886), .ZN(n_0_81_24));
   INV_X1 i_0_81_49 (.A(n_0_81_24), .ZN(n_0_1983));
   AOI222_X1 i_0_81_50 (.A1(n_0_1958), .A2(n_0_1950), .B1(n_0_1959), .B2(
      n_0_1918), .C1(n_0_1957), .C2(n_0_1887), .ZN(n_0_81_25));
   INV_X1 i_0_81_51 (.A(n_0_81_25), .ZN(n_0_1984));
   AOI222_X1 i_0_81_52 (.A1(n_0_1958), .A2(n_0_1951), .B1(n_0_1959), .B2(
      n_0_1919), .C1(n_0_1957), .C2(n_0_1888), .ZN(n_0_81_26));
   INV_X1 i_0_81_53 (.A(n_0_81_26), .ZN(n_0_1985));
   AOI222_X1 i_0_81_54 (.A1(n_0_1958), .A2(n_0_1952), .B1(n_0_1959), .B2(
      n_0_1920), .C1(n_0_1957), .C2(n_0_1889), .ZN(n_0_81_27));
   INV_X1 i_0_81_55 (.A(n_0_81_27), .ZN(n_0_1986));
   AOI222_X1 i_0_81_56 (.A1(n_0_1958), .A2(n_0_1953), .B1(n_0_1959), .B2(
      n_0_1921), .C1(n_0_1957), .C2(n_0_1890), .ZN(n_0_81_28));
   INV_X1 i_0_81_57 (.A(n_0_81_28), .ZN(n_0_1987));
   AOI222_X1 i_0_81_58 (.A1(n_0_1958), .A2(n_0_1954), .B1(n_0_1959), .B2(
      n_0_1922), .C1(n_0_1957), .C2(n_0_1891), .ZN(n_0_81_29));
   INV_X1 i_0_81_59 (.A(n_0_81_29), .ZN(n_0_1988));
   AND2_X1 i_0_81_60 (.A1(n_0_1957), .A2(n_0_1892), .ZN(n_0_81_30));
   AOI221_X1 i_0_81_61 (.A(n_0_81_30), .B1(n_0_1958), .B2(n_0_1955), .C1(
      n_0_1959), .C2(n_0_1923), .ZN(n_0_81_31));
   INV_X1 i_0_81_62 (.A(n_0_81_31), .ZN(n_0_1989));
   AOI221_X1 i_0_81_63 (.A(n_0_81_30), .B1(n_0_1958), .B2(n_0_1956), .C1(
      n_0_1959), .C2(n_0_1924), .ZN(n_0_81_32));
   INV_X1 i_0_81_64 (.A(n_0_81_32), .ZN(n_0_1990));
   datapath__0_80 i_0_82 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_41, 
      n_0_1990, n_0_1989, n_0_1988, n_0_1987, n_0_1986, n_0_1985, n_0_1984, 
      n_0_1983, n_0_1982, n_0_1981, n_0_1980, n_0_1979, n_0_1978, n_0_1977, 
      n_0_1976, n_0_1975, n_0_1974, n_0_1973, n_0_1972, n_0_1971, n_0_1970, 
      n_0_1969, n_0_1968, n_0_1967, n_0_1966, n_0_1965, n_0_1964, n_0_1963, 
      n_0_1962, n_0_1961, n_0_1960}), .p_2({n_0_2022, n_0_2021, n_0_2020, 
      n_0_2019, n_0_2018, n_0_2017, n_0_2016, n_0_2015, n_0_2014, n_0_2013, 
      n_0_2012, n_0_2011, n_0_2010, n_0_2009, n_0_2008, n_0_2007, n_0_2006, 
      n_0_2005, n_0_2004, n_0_2003, n_0_2002, n_0_2001, n_0_2000, n_0_1999, 
      n_0_1998, n_0_1997, n_0_1996, n_0_1995, n_0_1994, n_0_1993, n_0_1992, 
      n_0_1991}));
   datapath__0_81 i_0_83 (.multiplicand2(multiplicand2), .p_0({uc_42, n_0_1990, 
      n_0_1989, n_0_1988, n_0_1987, n_0_1986, n_0_1985, n_0_1984, n_0_1983, 
      n_0_1982, n_0_1981, n_0_1980, n_0_1979, n_0_1978, n_0_1977, n_0_1976, 
      n_0_1975, n_0_1974, n_0_1973, n_0_1972, n_0_1971, n_0_1970, n_0_1969, 
      n_0_1968, n_0_1967, n_0_1966, n_0_1965, n_0_1964, n_0_1963, n_0_1962, 
      n_0_1961, n_0_1960}), .p_1({n_0_2054, n_0_2053, n_0_2052, n_0_2051, 
      n_0_2050, n_0_2049, n_0_2048, n_0_2047, n_0_2046, n_0_2045, n_0_2044, 
      n_0_2043, n_0_2042, n_0_2041, n_0_2040, n_0_2039, n_0_2038, n_0_2037, 
      n_0_2036, n_0_2035, n_0_2034, n_0_2033, n_0_2032, n_0_2031, n_0_2030, 
      n_0_2029, n_0_2028, n_0_2027, n_0_2026, n_0_2025, n_0_2024, n_0_2023}));
   INV_X1 i_0_84_0 (.A(multiplier2[21]), .ZN(n_0_84_0));
   AND2_X1 i_0_84_1 (.A1(n_0_84_0), .A2(multiplier2[20]), .ZN(n_0_2056));
   NOR2_X1 i_0_84_2 (.A1(n_0_84_0), .A2(multiplier2[20]), .ZN(n_0_2057));
   NOR2_X1 i_0_84_3 (.A1(n_0_2056), .A2(n_0_2057), .ZN(n_0_2055));
   AOI222_X1 i_0_85_0 (.A1(n_0_2023), .A2(n_0_2056), .B1(n_0_1991), .B2(n_0_2057), 
      .C1(n_0_1960), .C2(n_0_2055), .ZN(n_0_85_0));
   INV_X1 i_0_85_1 (.A(n_0_85_0), .ZN(product[21]));
   AOI222_X1 i_0_85_2 (.A1(n_0_2056), .A2(n_0_2024), .B1(n_0_2057), .B2(n_0_1992), 
      .C1(n_0_2055), .C2(n_0_1961), .ZN(n_0_85_1));
   INV_X1 i_0_85_3 (.A(n_0_85_1), .ZN(n_0_2058));
   AOI222_X1 i_0_85_4 (.A1(n_0_2056), .A2(n_0_2025), .B1(n_0_2057), .B2(n_0_1993), 
      .C1(n_0_2055), .C2(n_0_1962), .ZN(n_0_85_2));
   INV_X1 i_0_85_5 (.A(n_0_85_2), .ZN(n_0_2059));
   AOI222_X1 i_0_85_6 (.A1(n_0_2056), .A2(n_0_2026), .B1(n_0_2057), .B2(n_0_1994), 
      .C1(n_0_2055), .C2(n_0_1963), .ZN(n_0_85_3));
   INV_X1 i_0_85_7 (.A(n_0_85_3), .ZN(n_0_2060));
   AOI222_X1 i_0_85_8 (.A1(n_0_2056), .A2(n_0_2027), .B1(n_0_2057), .B2(n_0_1995), 
      .C1(n_0_2055), .C2(n_0_1964), .ZN(n_0_85_4));
   INV_X1 i_0_85_9 (.A(n_0_85_4), .ZN(n_0_2061));
   AOI222_X1 i_0_85_10 (.A1(n_0_2056), .A2(n_0_2028), .B1(n_0_2057), .B2(
      n_0_1996), .C1(n_0_2055), .C2(n_0_1965), .ZN(n_0_85_5));
   INV_X1 i_0_85_11 (.A(n_0_85_5), .ZN(n_0_2062));
   AOI222_X1 i_0_85_12 (.A1(n_0_2056), .A2(n_0_2029), .B1(n_0_2057), .B2(
      n_0_1997), .C1(n_0_2055), .C2(n_0_1966), .ZN(n_0_85_6));
   INV_X1 i_0_85_13 (.A(n_0_85_6), .ZN(n_0_2063));
   AOI222_X1 i_0_85_14 (.A1(n_0_2056), .A2(n_0_2030), .B1(n_0_2057), .B2(
      n_0_1998), .C1(n_0_2055), .C2(n_0_1967), .ZN(n_0_85_7));
   INV_X1 i_0_85_15 (.A(n_0_85_7), .ZN(n_0_2064));
   AOI222_X1 i_0_85_16 (.A1(n_0_2056), .A2(n_0_2031), .B1(n_0_2057), .B2(
      n_0_1999), .C1(n_0_2055), .C2(n_0_1968), .ZN(n_0_85_8));
   INV_X1 i_0_85_17 (.A(n_0_85_8), .ZN(n_0_2065));
   AOI222_X1 i_0_85_18 (.A1(n_0_2056), .A2(n_0_2032), .B1(n_0_2057), .B2(
      n_0_2000), .C1(n_0_2055), .C2(n_0_1969), .ZN(n_0_85_9));
   INV_X1 i_0_85_19 (.A(n_0_85_9), .ZN(n_0_2066));
   AOI222_X1 i_0_85_20 (.A1(n_0_2056), .A2(n_0_2033), .B1(n_0_2057), .B2(
      n_0_2001), .C1(n_0_2055), .C2(n_0_1970), .ZN(n_0_85_10));
   INV_X1 i_0_85_21 (.A(n_0_85_10), .ZN(n_0_2067));
   AOI222_X1 i_0_85_22 (.A1(n_0_2056), .A2(n_0_2034), .B1(n_0_2057), .B2(
      n_0_2002), .C1(n_0_2055), .C2(n_0_1971), .ZN(n_0_85_11));
   INV_X1 i_0_85_23 (.A(n_0_85_11), .ZN(n_0_2068));
   AOI222_X1 i_0_85_24 (.A1(n_0_2056), .A2(n_0_2035), .B1(n_0_2057), .B2(
      n_0_2003), .C1(n_0_2055), .C2(n_0_1972), .ZN(n_0_85_12));
   INV_X1 i_0_85_25 (.A(n_0_85_12), .ZN(n_0_2069));
   AOI222_X1 i_0_85_26 (.A1(n_0_2056), .A2(n_0_2036), .B1(n_0_2057), .B2(
      n_0_2004), .C1(n_0_2055), .C2(n_0_1973), .ZN(n_0_85_13));
   INV_X1 i_0_85_27 (.A(n_0_85_13), .ZN(n_0_2070));
   AOI222_X1 i_0_85_28 (.A1(n_0_2056), .A2(n_0_2037), .B1(n_0_2057), .B2(
      n_0_2005), .C1(n_0_2055), .C2(n_0_1974), .ZN(n_0_85_14));
   INV_X1 i_0_85_29 (.A(n_0_85_14), .ZN(n_0_2071));
   AOI222_X1 i_0_85_30 (.A1(n_0_2056), .A2(n_0_2038), .B1(n_0_2057), .B2(
      n_0_2006), .C1(n_0_2055), .C2(n_0_1975), .ZN(n_0_85_15));
   INV_X1 i_0_85_31 (.A(n_0_85_15), .ZN(n_0_2072));
   AOI222_X1 i_0_85_32 (.A1(n_0_2056), .A2(n_0_2039), .B1(n_0_2057), .B2(
      n_0_2007), .C1(n_0_2055), .C2(n_0_1976), .ZN(n_0_85_16));
   INV_X1 i_0_85_33 (.A(n_0_85_16), .ZN(n_0_2073));
   AOI222_X1 i_0_85_34 (.A1(n_0_2056), .A2(n_0_2040), .B1(n_0_2057), .B2(
      n_0_2008), .C1(n_0_2055), .C2(n_0_1977), .ZN(n_0_85_17));
   INV_X1 i_0_85_35 (.A(n_0_85_17), .ZN(n_0_2074));
   AOI222_X1 i_0_85_36 (.A1(n_0_2056), .A2(n_0_2041), .B1(n_0_2057), .B2(
      n_0_2009), .C1(n_0_2055), .C2(n_0_1978), .ZN(n_0_85_18));
   INV_X1 i_0_85_37 (.A(n_0_85_18), .ZN(n_0_2075));
   AOI222_X1 i_0_85_38 (.A1(n_0_2056), .A2(n_0_2042), .B1(n_0_2057), .B2(
      n_0_2010), .C1(n_0_2055), .C2(n_0_1979), .ZN(n_0_85_19));
   INV_X1 i_0_85_39 (.A(n_0_85_19), .ZN(n_0_2076));
   AOI222_X1 i_0_85_40 (.A1(n_0_2056), .A2(n_0_2043), .B1(n_0_2057), .B2(
      n_0_2011), .C1(n_0_2055), .C2(n_0_1980), .ZN(n_0_85_20));
   INV_X1 i_0_85_41 (.A(n_0_85_20), .ZN(n_0_2077));
   AOI222_X1 i_0_85_42 (.A1(n_0_2056), .A2(n_0_2044), .B1(n_0_2057), .B2(
      n_0_2012), .C1(n_0_2055), .C2(n_0_1981), .ZN(n_0_85_21));
   INV_X1 i_0_85_43 (.A(n_0_85_21), .ZN(n_0_2078));
   AOI222_X1 i_0_85_44 (.A1(n_0_2056), .A2(n_0_2045), .B1(n_0_2057), .B2(
      n_0_2013), .C1(n_0_2055), .C2(n_0_1982), .ZN(n_0_85_22));
   INV_X1 i_0_85_45 (.A(n_0_85_22), .ZN(n_0_2079));
   AOI222_X1 i_0_85_46 (.A1(n_0_2056), .A2(n_0_2046), .B1(n_0_2057), .B2(
      n_0_2014), .C1(n_0_2055), .C2(n_0_1983), .ZN(n_0_85_23));
   INV_X1 i_0_85_47 (.A(n_0_85_23), .ZN(n_0_2080));
   AOI222_X1 i_0_85_48 (.A1(n_0_2056), .A2(n_0_2047), .B1(n_0_2057), .B2(
      n_0_2015), .C1(n_0_2055), .C2(n_0_1984), .ZN(n_0_85_24));
   INV_X1 i_0_85_49 (.A(n_0_85_24), .ZN(n_0_2081));
   AOI222_X1 i_0_85_50 (.A1(n_0_2056), .A2(n_0_2048), .B1(n_0_2057), .B2(
      n_0_2016), .C1(n_0_2055), .C2(n_0_1985), .ZN(n_0_85_25));
   INV_X1 i_0_85_51 (.A(n_0_85_25), .ZN(n_0_2082));
   AOI222_X1 i_0_85_52 (.A1(n_0_2056), .A2(n_0_2049), .B1(n_0_2057), .B2(
      n_0_2017), .C1(n_0_2055), .C2(n_0_1986), .ZN(n_0_85_26));
   INV_X1 i_0_85_53 (.A(n_0_85_26), .ZN(n_0_2083));
   AOI222_X1 i_0_85_54 (.A1(n_0_2056), .A2(n_0_2050), .B1(n_0_2057), .B2(
      n_0_2018), .C1(n_0_2055), .C2(n_0_1987), .ZN(n_0_85_27));
   INV_X1 i_0_85_55 (.A(n_0_85_27), .ZN(n_0_2084));
   AOI222_X1 i_0_85_56 (.A1(n_0_2056), .A2(n_0_2051), .B1(n_0_2057), .B2(
      n_0_2019), .C1(n_0_2055), .C2(n_0_1988), .ZN(n_0_85_28));
   INV_X1 i_0_85_57 (.A(n_0_85_28), .ZN(n_0_2085));
   AOI222_X1 i_0_85_58 (.A1(n_0_2056), .A2(n_0_2052), .B1(n_0_2057), .B2(
      n_0_2020), .C1(n_0_2055), .C2(n_0_1989), .ZN(n_0_85_29));
   INV_X1 i_0_85_59 (.A(n_0_85_29), .ZN(n_0_2086));
   AND2_X1 i_0_85_60 (.A1(n_0_2055), .A2(n_0_1990), .ZN(n_0_85_30));
   AOI221_X1 i_0_85_61 (.A(n_0_85_30), .B1(n_0_2056), .B2(n_0_2053), .C1(
      n_0_2057), .C2(n_0_2021), .ZN(n_0_85_31));
   INV_X1 i_0_85_62 (.A(n_0_85_31), .ZN(n_0_2087));
   AOI221_X1 i_0_85_63 (.A(n_0_85_30), .B1(n_0_2056), .B2(n_0_2054), .C1(
      n_0_2057), .C2(n_0_2022), .ZN(n_0_85_32));
   INV_X1 i_0_85_64 (.A(n_0_85_32), .ZN(n_0_2088));
   datapath__0_84 i_0_86 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_43, 
      n_0_2088, n_0_2087, n_0_2086, n_0_2085, n_0_2084, n_0_2083, n_0_2082, 
      n_0_2081, n_0_2080, n_0_2079, n_0_2078, n_0_2077, n_0_2076, n_0_2075, 
      n_0_2074, n_0_2073, n_0_2072, n_0_2071, n_0_2070, n_0_2069, n_0_2068, 
      n_0_2067, n_0_2066, n_0_2065, n_0_2064, n_0_2063, n_0_2062, n_0_2061, 
      n_0_2060, n_0_2059, n_0_2058}), .p_2({n_0_2120, n_0_2119, n_0_2118, 
      n_0_2117, n_0_2116, n_0_2115, n_0_2114, n_0_2113, n_0_2112, n_0_2111, 
      n_0_2110, n_0_2109, n_0_2108, n_0_2107, n_0_2106, n_0_2105, n_0_2104, 
      n_0_2103, n_0_2102, n_0_2101, n_0_2100, n_0_2099, n_0_2098, n_0_2097, 
      n_0_2096, n_0_2095, n_0_2094, n_0_2093, n_0_2092, n_0_2091, n_0_2090, 
      n_0_2089}));
   datapath__0_85 i_0_87 (.multiplicand2(multiplicand2), .p_0({uc_44, n_0_2088, 
      n_0_2087, n_0_2086, n_0_2085, n_0_2084, n_0_2083, n_0_2082, n_0_2081, 
      n_0_2080, n_0_2079, n_0_2078, n_0_2077, n_0_2076, n_0_2075, n_0_2074, 
      n_0_2073, n_0_2072, n_0_2071, n_0_2070, n_0_2069, n_0_2068, n_0_2067, 
      n_0_2066, n_0_2065, n_0_2064, n_0_2063, n_0_2062, n_0_2061, n_0_2060, 
      n_0_2059, n_0_2058}), .p_1({n_0_2152, n_0_2151, n_0_2150, n_0_2149, 
      n_0_2148, n_0_2147, n_0_2146, n_0_2145, n_0_2144, n_0_2143, n_0_2142, 
      n_0_2141, n_0_2140, n_0_2139, n_0_2138, n_0_2137, n_0_2136, n_0_2135, 
      n_0_2134, n_0_2133, n_0_2132, n_0_2131, n_0_2130, n_0_2129, n_0_2128, 
      n_0_2127, n_0_2126, n_0_2125, n_0_2124, n_0_2123, n_0_2122, n_0_2121}));
   INV_X1 i_0_88_0 (.A(multiplier2[22]), .ZN(n_0_88_0));
   AND2_X1 i_0_88_1 (.A1(n_0_88_0), .A2(multiplier2[21]), .ZN(n_0_2154));
   NOR2_X1 i_0_88_2 (.A1(n_0_88_0), .A2(multiplier2[21]), .ZN(n_0_2155));
   NOR2_X1 i_0_88_3 (.A1(n_0_2154), .A2(n_0_2155), .ZN(n_0_2153));
   AOI222_X1 i_0_89_0 (.A1(n_0_2121), .A2(n_0_2154), .B1(n_0_2089), .B2(n_0_2155), 
      .C1(n_0_2058), .C2(n_0_2153), .ZN(n_0_89_0));
   INV_X1 i_0_89_1 (.A(n_0_89_0), .ZN(product[22]));
   AOI222_X1 i_0_89_2 (.A1(n_0_2154), .A2(n_0_2122), .B1(n_0_2155), .B2(n_0_2090), 
      .C1(n_0_2153), .C2(n_0_2059), .ZN(n_0_89_1));
   INV_X1 i_0_89_3 (.A(n_0_89_1), .ZN(n_0_2156));
   AOI222_X1 i_0_89_4 (.A1(n_0_2154), .A2(n_0_2123), .B1(n_0_2155), .B2(n_0_2091), 
      .C1(n_0_2153), .C2(n_0_2060), .ZN(n_0_89_2));
   INV_X1 i_0_89_5 (.A(n_0_89_2), .ZN(n_0_2157));
   AOI222_X1 i_0_89_6 (.A1(n_0_2154), .A2(n_0_2124), .B1(n_0_2155), .B2(n_0_2092), 
      .C1(n_0_2153), .C2(n_0_2061), .ZN(n_0_89_3));
   INV_X1 i_0_89_7 (.A(n_0_89_3), .ZN(n_0_2158));
   AOI222_X1 i_0_89_8 (.A1(n_0_2154), .A2(n_0_2125), .B1(n_0_2155), .B2(n_0_2093), 
      .C1(n_0_2153), .C2(n_0_2062), .ZN(n_0_89_4));
   INV_X1 i_0_89_9 (.A(n_0_89_4), .ZN(n_0_2159));
   AOI222_X1 i_0_89_10 (.A1(n_0_2154), .A2(n_0_2126), .B1(n_0_2155), .B2(
      n_0_2094), .C1(n_0_2153), .C2(n_0_2063), .ZN(n_0_89_5));
   INV_X1 i_0_89_11 (.A(n_0_89_5), .ZN(n_0_2160));
   AOI222_X1 i_0_89_12 (.A1(n_0_2154), .A2(n_0_2127), .B1(n_0_2155), .B2(
      n_0_2095), .C1(n_0_2153), .C2(n_0_2064), .ZN(n_0_89_6));
   INV_X1 i_0_89_13 (.A(n_0_89_6), .ZN(n_0_2161));
   AOI222_X1 i_0_89_14 (.A1(n_0_2154), .A2(n_0_2128), .B1(n_0_2155), .B2(
      n_0_2096), .C1(n_0_2153), .C2(n_0_2065), .ZN(n_0_89_7));
   INV_X1 i_0_89_15 (.A(n_0_89_7), .ZN(n_0_2162));
   AOI222_X1 i_0_89_16 (.A1(n_0_2154), .A2(n_0_2129), .B1(n_0_2155), .B2(
      n_0_2097), .C1(n_0_2153), .C2(n_0_2066), .ZN(n_0_89_8));
   INV_X1 i_0_89_17 (.A(n_0_89_8), .ZN(n_0_2163));
   AOI222_X1 i_0_89_18 (.A1(n_0_2154), .A2(n_0_2130), .B1(n_0_2155), .B2(
      n_0_2098), .C1(n_0_2153), .C2(n_0_2067), .ZN(n_0_89_9));
   INV_X1 i_0_89_19 (.A(n_0_89_9), .ZN(n_0_2164));
   AOI222_X1 i_0_89_20 (.A1(n_0_2154), .A2(n_0_2131), .B1(n_0_2155), .B2(
      n_0_2099), .C1(n_0_2153), .C2(n_0_2068), .ZN(n_0_89_10));
   INV_X1 i_0_89_21 (.A(n_0_89_10), .ZN(n_0_2165));
   AOI222_X1 i_0_89_22 (.A1(n_0_2154), .A2(n_0_2132), .B1(n_0_2155), .B2(
      n_0_2100), .C1(n_0_2153), .C2(n_0_2069), .ZN(n_0_89_11));
   INV_X1 i_0_89_23 (.A(n_0_89_11), .ZN(n_0_2166));
   AOI222_X1 i_0_89_24 (.A1(n_0_2154), .A2(n_0_2133), .B1(n_0_2155), .B2(
      n_0_2101), .C1(n_0_2153), .C2(n_0_2070), .ZN(n_0_89_12));
   INV_X1 i_0_89_25 (.A(n_0_89_12), .ZN(n_0_2167));
   AOI222_X1 i_0_89_26 (.A1(n_0_2154), .A2(n_0_2134), .B1(n_0_2155), .B2(
      n_0_2102), .C1(n_0_2153), .C2(n_0_2071), .ZN(n_0_89_13));
   INV_X1 i_0_89_27 (.A(n_0_89_13), .ZN(n_0_2168));
   AOI222_X1 i_0_89_28 (.A1(n_0_2154), .A2(n_0_2135), .B1(n_0_2155), .B2(
      n_0_2103), .C1(n_0_2153), .C2(n_0_2072), .ZN(n_0_89_14));
   INV_X1 i_0_89_29 (.A(n_0_89_14), .ZN(n_0_2169));
   AOI222_X1 i_0_89_30 (.A1(n_0_2154), .A2(n_0_2136), .B1(n_0_2155), .B2(
      n_0_2104), .C1(n_0_2153), .C2(n_0_2073), .ZN(n_0_89_15));
   INV_X1 i_0_89_31 (.A(n_0_89_15), .ZN(n_0_2170));
   AOI222_X1 i_0_89_32 (.A1(n_0_2154), .A2(n_0_2137), .B1(n_0_2155), .B2(
      n_0_2105), .C1(n_0_2153), .C2(n_0_2074), .ZN(n_0_89_16));
   INV_X1 i_0_89_33 (.A(n_0_89_16), .ZN(n_0_2171));
   AOI222_X1 i_0_89_34 (.A1(n_0_2154), .A2(n_0_2138), .B1(n_0_2155), .B2(
      n_0_2106), .C1(n_0_2153), .C2(n_0_2075), .ZN(n_0_89_17));
   INV_X1 i_0_89_35 (.A(n_0_89_17), .ZN(n_0_2172));
   AOI222_X1 i_0_89_36 (.A1(n_0_2154), .A2(n_0_2139), .B1(n_0_2155), .B2(
      n_0_2107), .C1(n_0_2153), .C2(n_0_2076), .ZN(n_0_89_18));
   INV_X1 i_0_89_37 (.A(n_0_89_18), .ZN(n_0_2173));
   AOI222_X1 i_0_89_38 (.A1(n_0_2154), .A2(n_0_2140), .B1(n_0_2155), .B2(
      n_0_2108), .C1(n_0_2153), .C2(n_0_2077), .ZN(n_0_89_19));
   INV_X1 i_0_89_39 (.A(n_0_89_19), .ZN(n_0_2174));
   AOI222_X1 i_0_89_40 (.A1(n_0_2154), .A2(n_0_2141), .B1(n_0_2155), .B2(
      n_0_2109), .C1(n_0_2153), .C2(n_0_2078), .ZN(n_0_89_20));
   INV_X1 i_0_89_41 (.A(n_0_89_20), .ZN(n_0_2175));
   AOI222_X1 i_0_89_42 (.A1(n_0_2154), .A2(n_0_2142), .B1(n_0_2155), .B2(
      n_0_2110), .C1(n_0_2153), .C2(n_0_2079), .ZN(n_0_89_21));
   INV_X1 i_0_89_43 (.A(n_0_89_21), .ZN(n_0_2176));
   AOI222_X1 i_0_89_44 (.A1(n_0_2154), .A2(n_0_2143), .B1(n_0_2155), .B2(
      n_0_2111), .C1(n_0_2153), .C2(n_0_2080), .ZN(n_0_89_22));
   INV_X1 i_0_89_45 (.A(n_0_89_22), .ZN(n_0_2177));
   AOI222_X1 i_0_89_46 (.A1(n_0_2154), .A2(n_0_2144), .B1(n_0_2155), .B2(
      n_0_2112), .C1(n_0_2153), .C2(n_0_2081), .ZN(n_0_89_23));
   INV_X1 i_0_89_47 (.A(n_0_89_23), .ZN(n_0_2178));
   AOI222_X1 i_0_89_48 (.A1(n_0_2154), .A2(n_0_2145), .B1(n_0_2155), .B2(
      n_0_2113), .C1(n_0_2153), .C2(n_0_2082), .ZN(n_0_89_24));
   INV_X1 i_0_89_49 (.A(n_0_89_24), .ZN(n_0_2179));
   AOI222_X1 i_0_89_50 (.A1(n_0_2154), .A2(n_0_2146), .B1(n_0_2155), .B2(
      n_0_2114), .C1(n_0_2153), .C2(n_0_2083), .ZN(n_0_89_25));
   INV_X1 i_0_89_51 (.A(n_0_89_25), .ZN(n_0_2180));
   AOI222_X1 i_0_89_52 (.A1(n_0_2154), .A2(n_0_2147), .B1(n_0_2155), .B2(
      n_0_2115), .C1(n_0_2153), .C2(n_0_2084), .ZN(n_0_89_26));
   INV_X1 i_0_89_53 (.A(n_0_89_26), .ZN(n_0_2181));
   AOI222_X1 i_0_89_54 (.A1(n_0_2154), .A2(n_0_2148), .B1(n_0_2155), .B2(
      n_0_2116), .C1(n_0_2153), .C2(n_0_2085), .ZN(n_0_89_27));
   INV_X1 i_0_89_55 (.A(n_0_89_27), .ZN(n_0_2182));
   AOI222_X1 i_0_89_56 (.A1(n_0_2154), .A2(n_0_2149), .B1(n_0_2155), .B2(
      n_0_2117), .C1(n_0_2153), .C2(n_0_2086), .ZN(n_0_89_28));
   INV_X1 i_0_89_57 (.A(n_0_89_28), .ZN(n_0_2183));
   AOI222_X1 i_0_89_58 (.A1(n_0_2154), .A2(n_0_2150), .B1(n_0_2155), .B2(
      n_0_2118), .C1(n_0_2153), .C2(n_0_2087), .ZN(n_0_89_29));
   INV_X1 i_0_89_59 (.A(n_0_89_29), .ZN(n_0_2184));
   AND2_X1 i_0_89_60 (.A1(n_0_2153), .A2(n_0_2088), .ZN(n_0_89_30));
   AOI221_X1 i_0_89_61 (.A(n_0_89_30), .B1(n_0_2154), .B2(n_0_2151), .C1(
      n_0_2155), .C2(n_0_2119), .ZN(n_0_89_31));
   INV_X1 i_0_89_62 (.A(n_0_89_31), .ZN(n_0_2185));
   AOI221_X1 i_0_89_63 (.A(n_0_89_30), .B1(n_0_2154), .B2(n_0_2152), .C1(
      n_0_2155), .C2(n_0_2120), .ZN(n_0_89_32));
   INV_X1 i_0_89_64 (.A(n_0_89_32), .ZN(n_0_2186));
   datapath__0_88 i_0_90 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_45, 
      n_0_2186, n_0_2185, n_0_2184, n_0_2183, n_0_2182, n_0_2181, n_0_2180, 
      n_0_2179, n_0_2178, n_0_2177, n_0_2176, n_0_2175, n_0_2174, n_0_2173, 
      n_0_2172, n_0_2171, n_0_2170, n_0_2169, n_0_2168, n_0_2167, n_0_2166, 
      n_0_2165, n_0_2164, n_0_2163, n_0_2162, n_0_2161, n_0_2160, n_0_2159, 
      n_0_2158, n_0_2157, n_0_2156}), .p_2({n_0_2218, n_0_2217, n_0_2216, 
      n_0_2215, n_0_2214, n_0_2213, n_0_2212, n_0_2211, n_0_2210, n_0_2209, 
      n_0_2208, n_0_2207, n_0_2206, n_0_2205, n_0_2204, n_0_2203, n_0_2202, 
      n_0_2201, n_0_2200, n_0_2199, n_0_2198, n_0_2197, n_0_2196, n_0_2195, 
      n_0_2194, n_0_2193, n_0_2192, n_0_2191, n_0_2190, n_0_2189, n_0_2188, 
      n_0_2187}));
   datapath__0_89 i_0_91 (.multiplicand2(multiplicand2), .p_0({uc_46, n_0_2186, 
      n_0_2185, n_0_2184, n_0_2183, n_0_2182, n_0_2181, n_0_2180, n_0_2179, 
      n_0_2178, n_0_2177, n_0_2176, n_0_2175, n_0_2174, n_0_2173, n_0_2172, 
      n_0_2171, n_0_2170, n_0_2169, n_0_2168, n_0_2167, n_0_2166, n_0_2165, 
      n_0_2164, n_0_2163, n_0_2162, n_0_2161, n_0_2160, n_0_2159, n_0_2158, 
      n_0_2157, n_0_2156}), .p_1({n_0_2250, n_0_2249, n_0_2248, n_0_2247, 
      n_0_2246, n_0_2245, n_0_2244, n_0_2243, n_0_2242, n_0_2241, n_0_2240, 
      n_0_2239, n_0_2238, n_0_2237, n_0_2236, n_0_2235, n_0_2234, n_0_2233, 
      n_0_2232, n_0_2231, n_0_2230, n_0_2229, n_0_2228, n_0_2227, n_0_2226, 
      n_0_2225, n_0_2224, n_0_2223, n_0_2222, n_0_2221, n_0_2220, n_0_2219}));
   INV_X1 i_0_92_0 (.A(multiplier2[23]), .ZN(n_0_92_0));
   AND2_X1 i_0_92_1 (.A1(n_0_92_0), .A2(multiplier2[22]), .ZN(n_0_2252));
   NOR2_X1 i_0_92_2 (.A1(n_0_92_0), .A2(multiplier2[22]), .ZN(n_0_2253));
   NOR2_X1 i_0_92_3 (.A1(n_0_2252), .A2(n_0_2253), .ZN(n_0_2251));
   AOI222_X1 i_0_93_0 (.A1(n_0_2219), .A2(n_0_2252), .B1(n_0_2187), .B2(n_0_2253), 
      .C1(n_0_2156), .C2(n_0_2251), .ZN(n_0_93_0));
   INV_X1 i_0_93_1 (.A(n_0_93_0), .ZN(product[23]));
   AOI222_X1 i_0_93_2 (.A1(n_0_2252), .A2(n_0_2220), .B1(n_0_2253), .B2(n_0_2188), 
      .C1(n_0_2251), .C2(n_0_2157), .ZN(n_0_93_1));
   INV_X1 i_0_93_3 (.A(n_0_93_1), .ZN(n_0_2254));
   AOI222_X1 i_0_93_4 (.A1(n_0_2252), .A2(n_0_2221), .B1(n_0_2253), .B2(n_0_2189), 
      .C1(n_0_2251), .C2(n_0_2158), .ZN(n_0_93_2));
   INV_X1 i_0_93_5 (.A(n_0_93_2), .ZN(n_0_2255));
   AOI222_X1 i_0_93_6 (.A1(n_0_2252), .A2(n_0_2222), .B1(n_0_2253), .B2(n_0_2190), 
      .C1(n_0_2251), .C2(n_0_2159), .ZN(n_0_93_3));
   INV_X1 i_0_93_7 (.A(n_0_93_3), .ZN(n_0_2256));
   AOI222_X1 i_0_93_8 (.A1(n_0_2252), .A2(n_0_2223), .B1(n_0_2253), .B2(n_0_2191), 
      .C1(n_0_2251), .C2(n_0_2160), .ZN(n_0_93_4));
   INV_X1 i_0_93_9 (.A(n_0_93_4), .ZN(n_0_2257));
   AOI222_X1 i_0_93_10 (.A1(n_0_2252), .A2(n_0_2224), .B1(n_0_2253), .B2(
      n_0_2192), .C1(n_0_2251), .C2(n_0_2161), .ZN(n_0_93_5));
   INV_X1 i_0_93_11 (.A(n_0_93_5), .ZN(n_0_2258));
   AOI222_X1 i_0_93_12 (.A1(n_0_2252), .A2(n_0_2225), .B1(n_0_2253), .B2(
      n_0_2193), .C1(n_0_2251), .C2(n_0_2162), .ZN(n_0_93_6));
   INV_X1 i_0_93_13 (.A(n_0_93_6), .ZN(n_0_2259));
   AOI222_X1 i_0_93_14 (.A1(n_0_2252), .A2(n_0_2226), .B1(n_0_2253), .B2(
      n_0_2194), .C1(n_0_2251), .C2(n_0_2163), .ZN(n_0_93_7));
   INV_X1 i_0_93_15 (.A(n_0_93_7), .ZN(n_0_2260));
   AOI222_X1 i_0_93_16 (.A1(n_0_2252), .A2(n_0_2227), .B1(n_0_2253), .B2(
      n_0_2195), .C1(n_0_2251), .C2(n_0_2164), .ZN(n_0_93_8));
   INV_X1 i_0_93_17 (.A(n_0_93_8), .ZN(n_0_2261));
   AOI222_X1 i_0_93_18 (.A1(n_0_2252), .A2(n_0_2228), .B1(n_0_2253), .B2(
      n_0_2196), .C1(n_0_2251), .C2(n_0_2165), .ZN(n_0_93_9));
   INV_X1 i_0_93_19 (.A(n_0_93_9), .ZN(n_0_2262));
   AOI222_X1 i_0_93_20 (.A1(n_0_2252), .A2(n_0_2229), .B1(n_0_2253), .B2(
      n_0_2197), .C1(n_0_2251), .C2(n_0_2166), .ZN(n_0_93_10));
   INV_X1 i_0_93_21 (.A(n_0_93_10), .ZN(n_0_2263));
   AOI222_X1 i_0_93_22 (.A1(n_0_2252), .A2(n_0_2230), .B1(n_0_2253), .B2(
      n_0_2198), .C1(n_0_2251), .C2(n_0_2167), .ZN(n_0_93_11));
   INV_X1 i_0_93_23 (.A(n_0_93_11), .ZN(n_0_2264));
   AOI222_X1 i_0_93_24 (.A1(n_0_2252), .A2(n_0_2231), .B1(n_0_2253), .B2(
      n_0_2199), .C1(n_0_2251), .C2(n_0_2168), .ZN(n_0_93_12));
   INV_X1 i_0_93_25 (.A(n_0_93_12), .ZN(n_0_2265));
   AOI222_X1 i_0_93_26 (.A1(n_0_2252), .A2(n_0_2232), .B1(n_0_2253), .B2(
      n_0_2200), .C1(n_0_2251), .C2(n_0_2169), .ZN(n_0_93_13));
   INV_X1 i_0_93_27 (.A(n_0_93_13), .ZN(n_0_2266));
   AOI222_X1 i_0_93_28 (.A1(n_0_2252), .A2(n_0_2233), .B1(n_0_2253), .B2(
      n_0_2201), .C1(n_0_2251), .C2(n_0_2170), .ZN(n_0_93_14));
   INV_X1 i_0_93_29 (.A(n_0_93_14), .ZN(n_0_2267));
   AOI222_X1 i_0_93_30 (.A1(n_0_2252), .A2(n_0_2234), .B1(n_0_2253), .B2(
      n_0_2202), .C1(n_0_2251), .C2(n_0_2171), .ZN(n_0_93_15));
   INV_X1 i_0_93_31 (.A(n_0_93_15), .ZN(n_0_2268));
   AOI222_X1 i_0_93_32 (.A1(n_0_2252), .A2(n_0_2235), .B1(n_0_2253), .B2(
      n_0_2203), .C1(n_0_2251), .C2(n_0_2172), .ZN(n_0_93_16));
   INV_X1 i_0_93_33 (.A(n_0_93_16), .ZN(n_0_2269));
   AOI222_X1 i_0_93_34 (.A1(n_0_2252), .A2(n_0_2236), .B1(n_0_2253), .B2(
      n_0_2204), .C1(n_0_2251), .C2(n_0_2173), .ZN(n_0_93_17));
   INV_X1 i_0_93_35 (.A(n_0_93_17), .ZN(n_0_2270));
   AOI222_X1 i_0_93_36 (.A1(n_0_2252), .A2(n_0_2237), .B1(n_0_2253), .B2(
      n_0_2205), .C1(n_0_2251), .C2(n_0_2174), .ZN(n_0_93_18));
   INV_X1 i_0_93_37 (.A(n_0_93_18), .ZN(n_0_2271));
   AOI222_X1 i_0_93_38 (.A1(n_0_2252), .A2(n_0_2238), .B1(n_0_2253), .B2(
      n_0_2206), .C1(n_0_2251), .C2(n_0_2175), .ZN(n_0_93_19));
   INV_X1 i_0_93_39 (.A(n_0_93_19), .ZN(n_0_2272));
   AOI222_X1 i_0_93_40 (.A1(n_0_2252), .A2(n_0_2239), .B1(n_0_2253), .B2(
      n_0_2207), .C1(n_0_2251), .C2(n_0_2176), .ZN(n_0_93_20));
   INV_X1 i_0_93_41 (.A(n_0_93_20), .ZN(n_0_2273));
   AOI222_X1 i_0_93_42 (.A1(n_0_2252), .A2(n_0_2240), .B1(n_0_2253), .B2(
      n_0_2208), .C1(n_0_2251), .C2(n_0_2177), .ZN(n_0_93_21));
   INV_X1 i_0_93_43 (.A(n_0_93_21), .ZN(n_0_2274));
   AOI222_X1 i_0_93_44 (.A1(n_0_2252), .A2(n_0_2241), .B1(n_0_2253), .B2(
      n_0_2209), .C1(n_0_2251), .C2(n_0_2178), .ZN(n_0_93_22));
   INV_X1 i_0_93_45 (.A(n_0_93_22), .ZN(n_0_2275));
   AOI222_X1 i_0_93_46 (.A1(n_0_2252), .A2(n_0_2242), .B1(n_0_2253), .B2(
      n_0_2210), .C1(n_0_2251), .C2(n_0_2179), .ZN(n_0_93_23));
   INV_X1 i_0_93_47 (.A(n_0_93_23), .ZN(n_0_2276));
   AOI222_X1 i_0_93_48 (.A1(n_0_2252), .A2(n_0_2243), .B1(n_0_2253), .B2(
      n_0_2211), .C1(n_0_2251), .C2(n_0_2180), .ZN(n_0_93_24));
   INV_X1 i_0_93_49 (.A(n_0_93_24), .ZN(n_0_2277));
   AOI222_X1 i_0_93_50 (.A1(n_0_2252), .A2(n_0_2244), .B1(n_0_2253), .B2(
      n_0_2212), .C1(n_0_2251), .C2(n_0_2181), .ZN(n_0_93_25));
   INV_X1 i_0_93_51 (.A(n_0_93_25), .ZN(n_0_2278));
   AOI222_X1 i_0_93_52 (.A1(n_0_2252), .A2(n_0_2245), .B1(n_0_2253), .B2(
      n_0_2213), .C1(n_0_2251), .C2(n_0_2182), .ZN(n_0_93_26));
   INV_X1 i_0_93_53 (.A(n_0_93_26), .ZN(n_0_2279));
   AOI222_X1 i_0_93_54 (.A1(n_0_2252), .A2(n_0_2246), .B1(n_0_2253), .B2(
      n_0_2214), .C1(n_0_2251), .C2(n_0_2183), .ZN(n_0_93_27));
   INV_X1 i_0_93_55 (.A(n_0_93_27), .ZN(n_0_2280));
   AOI222_X1 i_0_93_56 (.A1(n_0_2252), .A2(n_0_2247), .B1(n_0_2253), .B2(
      n_0_2215), .C1(n_0_2251), .C2(n_0_2184), .ZN(n_0_93_28));
   INV_X1 i_0_93_57 (.A(n_0_93_28), .ZN(n_0_2281));
   AOI222_X1 i_0_93_58 (.A1(n_0_2252), .A2(n_0_2248), .B1(n_0_2253), .B2(
      n_0_2216), .C1(n_0_2251), .C2(n_0_2185), .ZN(n_0_93_29));
   INV_X1 i_0_93_59 (.A(n_0_93_29), .ZN(n_0_2282));
   AND2_X1 i_0_93_60 (.A1(n_0_2251), .A2(n_0_2186), .ZN(n_0_93_30));
   AOI221_X1 i_0_93_61 (.A(n_0_93_30), .B1(n_0_2252), .B2(n_0_2249), .C1(
      n_0_2253), .C2(n_0_2217), .ZN(n_0_93_31));
   INV_X1 i_0_93_62 (.A(n_0_93_31), .ZN(n_0_2283));
   AOI221_X1 i_0_93_63 (.A(n_0_93_30), .B1(n_0_2252), .B2(n_0_2250), .C1(
      n_0_2253), .C2(n_0_2218), .ZN(n_0_93_32));
   INV_X1 i_0_93_64 (.A(n_0_93_32), .ZN(n_0_2284));
   datapath__0_92 i_0_94 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_47, 
      n_0_2284, n_0_2283, n_0_2282, n_0_2281, n_0_2280, n_0_2279, n_0_2278, 
      n_0_2277, n_0_2276, n_0_2275, n_0_2274, n_0_2273, n_0_2272, n_0_2271, 
      n_0_2270, n_0_2269, n_0_2268, n_0_2267, n_0_2266, n_0_2265, n_0_2264, 
      n_0_2263, n_0_2262, n_0_2261, n_0_2260, n_0_2259, n_0_2258, n_0_2257, 
      n_0_2256, n_0_2255, n_0_2254}), .p_2({n_0_2316, n_0_2315, n_0_2314, 
      n_0_2313, n_0_2312, n_0_2311, n_0_2310, n_0_2309, n_0_2308, n_0_2307, 
      n_0_2306, n_0_2305, n_0_2304, n_0_2303, n_0_2302, n_0_2301, n_0_2300, 
      n_0_2299, n_0_2298, n_0_2297, n_0_2296, n_0_2295, n_0_2294, n_0_2293, 
      n_0_2292, n_0_2291, n_0_2290, n_0_2289, n_0_2288, n_0_2287, n_0_2286, 
      n_0_2285}));
   datapath__0_93 i_0_95 (.multiplicand2(multiplicand2), .p_0({uc_48, n_0_2284, 
      n_0_2283, n_0_2282, n_0_2281, n_0_2280, n_0_2279, n_0_2278, n_0_2277, 
      n_0_2276, n_0_2275, n_0_2274, n_0_2273, n_0_2272, n_0_2271, n_0_2270, 
      n_0_2269, n_0_2268, n_0_2267, n_0_2266, n_0_2265, n_0_2264, n_0_2263, 
      n_0_2262, n_0_2261, n_0_2260, n_0_2259, n_0_2258, n_0_2257, n_0_2256, 
      n_0_2255, n_0_2254}), .p_1({n_0_2348, n_0_2347, n_0_2346, n_0_2345, 
      n_0_2344, n_0_2343, n_0_2342, n_0_2341, n_0_2340, n_0_2339, n_0_2338, 
      n_0_2337, n_0_2336, n_0_2335, n_0_2334, n_0_2333, n_0_2332, n_0_2331, 
      n_0_2330, n_0_2329, n_0_2328, n_0_2327, n_0_2326, n_0_2325, n_0_2324, 
      n_0_2323, n_0_2322, n_0_2321, n_0_2320, n_0_2319, n_0_2318, n_0_2317}));
   INV_X1 i_0_96_0 (.A(multiplier2[24]), .ZN(n_0_96_0));
   AND2_X1 i_0_96_1 (.A1(n_0_96_0), .A2(multiplier2[23]), .ZN(n_0_2350));
   NOR2_X1 i_0_96_2 (.A1(n_0_96_0), .A2(multiplier2[23]), .ZN(n_0_2351));
   NOR2_X1 i_0_96_3 (.A1(n_0_2350), .A2(n_0_2351), .ZN(n_0_2349));
   AOI222_X1 i_0_97_0 (.A1(n_0_2317), .A2(n_0_2350), .B1(n_0_2285), .B2(n_0_2351), 
      .C1(n_0_2254), .C2(n_0_2349), .ZN(n_0_97_0));
   INV_X1 i_0_97_1 (.A(n_0_97_0), .ZN(product[24]));
   AOI222_X1 i_0_97_2 (.A1(n_0_2350), .A2(n_0_2318), .B1(n_0_2351), .B2(n_0_2286), 
      .C1(n_0_2349), .C2(n_0_2255), .ZN(n_0_97_1));
   INV_X1 i_0_97_3 (.A(n_0_97_1), .ZN(n_0_2352));
   AOI222_X1 i_0_97_4 (.A1(n_0_2350), .A2(n_0_2319), .B1(n_0_2351), .B2(n_0_2287), 
      .C1(n_0_2349), .C2(n_0_2256), .ZN(n_0_97_2));
   INV_X1 i_0_97_5 (.A(n_0_97_2), .ZN(n_0_2353));
   AOI222_X1 i_0_97_6 (.A1(n_0_2350), .A2(n_0_2320), .B1(n_0_2351), .B2(n_0_2288), 
      .C1(n_0_2349), .C2(n_0_2257), .ZN(n_0_97_3));
   INV_X1 i_0_97_7 (.A(n_0_97_3), .ZN(n_0_2354));
   AOI222_X1 i_0_97_8 (.A1(n_0_2350), .A2(n_0_2321), .B1(n_0_2351), .B2(n_0_2289), 
      .C1(n_0_2349), .C2(n_0_2258), .ZN(n_0_97_4));
   INV_X1 i_0_97_9 (.A(n_0_97_4), .ZN(n_0_2355));
   AOI222_X1 i_0_97_10 (.A1(n_0_2350), .A2(n_0_2322), .B1(n_0_2351), .B2(
      n_0_2290), .C1(n_0_2349), .C2(n_0_2259), .ZN(n_0_97_5));
   INV_X1 i_0_97_11 (.A(n_0_97_5), .ZN(n_0_2356));
   AOI222_X1 i_0_97_12 (.A1(n_0_2350), .A2(n_0_2323), .B1(n_0_2351), .B2(
      n_0_2291), .C1(n_0_2349), .C2(n_0_2260), .ZN(n_0_97_6));
   INV_X1 i_0_97_13 (.A(n_0_97_6), .ZN(n_0_2357));
   AOI222_X1 i_0_97_14 (.A1(n_0_2350), .A2(n_0_2324), .B1(n_0_2351), .B2(
      n_0_2292), .C1(n_0_2349), .C2(n_0_2261), .ZN(n_0_97_7));
   INV_X1 i_0_97_15 (.A(n_0_97_7), .ZN(n_0_2358));
   AOI222_X1 i_0_97_16 (.A1(n_0_2350), .A2(n_0_2325), .B1(n_0_2351), .B2(
      n_0_2293), .C1(n_0_2349), .C2(n_0_2262), .ZN(n_0_97_8));
   INV_X1 i_0_97_17 (.A(n_0_97_8), .ZN(n_0_2359));
   AOI222_X1 i_0_97_18 (.A1(n_0_2350), .A2(n_0_2326), .B1(n_0_2351), .B2(
      n_0_2294), .C1(n_0_2349), .C2(n_0_2263), .ZN(n_0_97_9));
   INV_X1 i_0_97_19 (.A(n_0_97_9), .ZN(n_0_2360));
   AOI222_X1 i_0_97_20 (.A1(n_0_2350), .A2(n_0_2327), .B1(n_0_2351), .B2(
      n_0_2295), .C1(n_0_2349), .C2(n_0_2264), .ZN(n_0_97_10));
   INV_X1 i_0_97_21 (.A(n_0_97_10), .ZN(n_0_2361));
   AOI222_X1 i_0_97_22 (.A1(n_0_2350), .A2(n_0_2328), .B1(n_0_2351), .B2(
      n_0_2296), .C1(n_0_2349), .C2(n_0_2265), .ZN(n_0_97_11));
   INV_X1 i_0_97_23 (.A(n_0_97_11), .ZN(n_0_2362));
   AOI222_X1 i_0_97_24 (.A1(n_0_2350), .A2(n_0_2329), .B1(n_0_2351), .B2(
      n_0_2297), .C1(n_0_2349), .C2(n_0_2266), .ZN(n_0_97_12));
   INV_X1 i_0_97_25 (.A(n_0_97_12), .ZN(n_0_2363));
   AOI222_X1 i_0_97_26 (.A1(n_0_2350), .A2(n_0_2330), .B1(n_0_2351), .B2(
      n_0_2298), .C1(n_0_2349), .C2(n_0_2267), .ZN(n_0_97_13));
   INV_X1 i_0_97_27 (.A(n_0_97_13), .ZN(n_0_2364));
   AOI222_X1 i_0_97_28 (.A1(n_0_2350), .A2(n_0_2331), .B1(n_0_2351), .B2(
      n_0_2299), .C1(n_0_2349), .C2(n_0_2268), .ZN(n_0_97_14));
   INV_X1 i_0_97_29 (.A(n_0_97_14), .ZN(n_0_2365));
   AOI222_X1 i_0_97_30 (.A1(n_0_2350), .A2(n_0_2332), .B1(n_0_2351), .B2(
      n_0_2300), .C1(n_0_2349), .C2(n_0_2269), .ZN(n_0_97_15));
   INV_X1 i_0_97_31 (.A(n_0_97_15), .ZN(n_0_2366));
   AOI222_X1 i_0_97_32 (.A1(n_0_2350), .A2(n_0_2333), .B1(n_0_2351), .B2(
      n_0_2301), .C1(n_0_2349), .C2(n_0_2270), .ZN(n_0_97_16));
   INV_X1 i_0_97_33 (.A(n_0_97_16), .ZN(n_0_2367));
   AOI222_X1 i_0_97_34 (.A1(n_0_2350), .A2(n_0_2334), .B1(n_0_2351), .B2(
      n_0_2302), .C1(n_0_2349), .C2(n_0_2271), .ZN(n_0_97_17));
   INV_X1 i_0_97_35 (.A(n_0_97_17), .ZN(n_0_2368));
   AOI222_X1 i_0_97_36 (.A1(n_0_2350), .A2(n_0_2335), .B1(n_0_2351), .B2(
      n_0_2303), .C1(n_0_2349), .C2(n_0_2272), .ZN(n_0_97_18));
   INV_X1 i_0_97_37 (.A(n_0_97_18), .ZN(n_0_2369));
   AOI222_X1 i_0_97_38 (.A1(n_0_2350), .A2(n_0_2336), .B1(n_0_2351), .B2(
      n_0_2304), .C1(n_0_2349), .C2(n_0_2273), .ZN(n_0_97_19));
   INV_X1 i_0_97_39 (.A(n_0_97_19), .ZN(n_0_2370));
   AOI222_X1 i_0_97_40 (.A1(n_0_2350), .A2(n_0_2337), .B1(n_0_2351), .B2(
      n_0_2305), .C1(n_0_2349), .C2(n_0_2274), .ZN(n_0_97_20));
   INV_X1 i_0_97_41 (.A(n_0_97_20), .ZN(n_0_2371));
   AOI222_X1 i_0_97_42 (.A1(n_0_2350), .A2(n_0_2338), .B1(n_0_2351), .B2(
      n_0_2306), .C1(n_0_2349), .C2(n_0_2275), .ZN(n_0_97_21));
   INV_X1 i_0_97_43 (.A(n_0_97_21), .ZN(n_0_2372));
   AOI222_X1 i_0_97_44 (.A1(n_0_2350), .A2(n_0_2339), .B1(n_0_2351), .B2(
      n_0_2307), .C1(n_0_2349), .C2(n_0_2276), .ZN(n_0_97_22));
   INV_X1 i_0_97_45 (.A(n_0_97_22), .ZN(n_0_2373));
   AOI222_X1 i_0_97_46 (.A1(n_0_2350), .A2(n_0_2340), .B1(n_0_2351), .B2(
      n_0_2308), .C1(n_0_2349), .C2(n_0_2277), .ZN(n_0_97_23));
   INV_X1 i_0_97_47 (.A(n_0_97_23), .ZN(n_0_2374));
   AOI222_X1 i_0_97_48 (.A1(n_0_2350), .A2(n_0_2341), .B1(n_0_2351), .B2(
      n_0_2309), .C1(n_0_2349), .C2(n_0_2278), .ZN(n_0_97_24));
   INV_X1 i_0_97_49 (.A(n_0_97_24), .ZN(n_0_2375));
   AOI222_X1 i_0_97_50 (.A1(n_0_2350), .A2(n_0_2342), .B1(n_0_2351), .B2(
      n_0_2310), .C1(n_0_2349), .C2(n_0_2279), .ZN(n_0_97_25));
   INV_X1 i_0_97_51 (.A(n_0_97_25), .ZN(n_0_2376));
   AOI222_X1 i_0_97_52 (.A1(n_0_2350), .A2(n_0_2343), .B1(n_0_2351), .B2(
      n_0_2311), .C1(n_0_2349), .C2(n_0_2280), .ZN(n_0_97_26));
   INV_X1 i_0_97_53 (.A(n_0_97_26), .ZN(n_0_2377));
   AOI222_X1 i_0_97_54 (.A1(n_0_2350), .A2(n_0_2344), .B1(n_0_2351), .B2(
      n_0_2312), .C1(n_0_2349), .C2(n_0_2281), .ZN(n_0_97_27));
   INV_X1 i_0_97_55 (.A(n_0_97_27), .ZN(n_0_2378));
   AOI222_X1 i_0_97_56 (.A1(n_0_2350), .A2(n_0_2345), .B1(n_0_2351), .B2(
      n_0_2313), .C1(n_0_2349), .C2(n_0_2282), .ZN(n_0_97_28));
   INV_X1 i_0_97_57 (.A(n_0_97_28), .ZN(n_0_2379));
   AOI222_X1 i_0_97_58 (.A1(n_0_2350), .A2(n_0_2346), .B1(n_0_2351), .B2(
      n_0_2314), .C1(n_0_2349), .C2(n_0_2283), .ZN(n_0_97_29));
   INV_X1 i_0_97_59 (.A(n_0_97_29), .ZN(n_0_2380));
   AND2_X1 i_0_97_60 (.A1(n_0_2349), .A2(n_0_2284), .ZN(n_0_97_30));
   AOI221_X1 i_0_97_61 (.A(n_0_97_30), .B1(n_0_2350), .B2(n_0_2347), .C1(
      n_0_2351), .C2(n_0_2315), .ZN(n_0_97_31));
   INV_X1 i_0_97_62 (.A(n_0_97_31), .ZN(n_0_2381));
   AOI221_X1 i_0_97_63 (.A(n_0_97_30), .B1(n_0_2350), .B2(n_0_2348), .C1(
      n_0_2351), .C2(n_0_2316), .ZN(n_0_97_32));
   INV_X1 i_0_97_64 (.A(n_0_97_32), .ZN(n_0_2382));
   datapath__0_96 i_0_98 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_49, 
      n_0_2382, n_0_2381, n_0_2380, n_0_2379, n_0_2378, n_0_2377, n_0_2376, 
      n_0_2375, n_0_2374, n_0_2373, n_0_2372, n_0_2371, n_0_2370, n_0_2369, 
      n_0_2368, n_0_2367, n_0_2366, n_0_2365, n_0_2364, n_0_2363, n_0_2362, 
      n_0_2361, n_0_2360, n_0_2359, n_0_2358, n_0_2357, n_0_2356, n_0_2355, 
      n_0_2354, n_0_2353, n_0_2352}), .p_2({n_0_2414, n_0_2413, n_0_2412, 
      n_0_2411, n_0_2410, n_0_2409, n_0_2408, n_0_2407, n_0_2406, n_0_2405, 
      n_0_2404, n_0_2403, n_0_2402, n_0_2401, n_0_2400, n_0_2399, n_0_2398, 
      n_0_2397, n_0_2396, n_0_2395, n_0_2394, n_0_2393, n_0_2392, n_0_2391, 
      n_0_2390, n_0_2389, n_0_2388, n_0_2387, n_0_2386, n_0_2385, n_0_2384, 
      n_0_2383}));
   datapath__0_97 i_0_99 (.multiplicand2(multiplicand2), .p_0({uc_50, n_0_2382, 
      n_0_2381, n_0_2380, n_0_2379, n_0_2378, n_0_2377, n_0_2376, n_0_2375, 
      n_0_2374, n_0_2373, n_0_2372, n_0_2371, n_0_2370, n_0_2369, n_0_2368, 
      n_0_2367, n_0_2366, n_0_2365, n_0_2364, n_0_2363, n_0_2362, n_0_2361, 
      n_0_2360, n_0_2359, n_0_2358, n_0_2357, n_0_2356, n_0_2355, n_0_2354, 
      n_0_2353, n_0_2352}), .p_1({n_0_2446, n_0_2445, n_0_2444, n_0_2443, 
      n_0_2442, n_0_2441, n_0_2440, n_0_2439, n_0_2438, n_0_2437, n_0_2436, 
      n_0_2435, n_0_2434, n_0_2433, n_0_2432, n_0_2431, n_0_2430, n_0_2429, 
      n_0_2428, n_0_2427, n_0_2426, n_0_2425, n_0_2424, n_0_2423, n_0_2422, 
      n_0_2421, n_0_2420, n_0_2419, n_0_2418, n_0_2417, n_0_2416, n_0_2415}));
   INV_X1 i_0_100_0 (.A(multiplier2[25]), .ZN(n_0_100_0));
   AND2_X1 i_0_100_1 (.A1(n_0_100_0), .A2(multiplier2[24]), .ZN(n_0_2448));
   NOR2_X1 i_0_100_2 (.A1(n_0_100_0), .A2(multiplier2[24]), .ZN(n_0_2449));
   NOR2_X1 i_0_100_3 (.A1(n_0_2448), .A2(n_0_2449), .ZN(n_0_2447));
   AOI222_X1 i_0_101_0 (.A1(n_0_2415), .A2(n_0_2448), .B1(n_0_2383), .B2(
      n_0_2449), .C1(n_0_2352), .C2(n_0_2447), .ZN(n_0_101_0));
   INV_X1 i_0_101_1 (.A(n_0_101_0), .ZN(product[25]));
   AOI222_X1 i_0_101_2 (.A1(n_0_2448), .A2(n_0_2416), .B1(n_0_2449), .B2(
      n_0_2384), .C1(n_0_2447), .C2(n_0_2353), .ZN(n_0_101_1));
   INV_X1 i_0_101_3 (.A(n_0_101_1), .ZN(n_0_2450));
   AOI222_X1 i_0_101_4 (.A1(n_0_2448), .A2(n_0_2417), .B1(n_0_2449), .B2(
      n_0_2385), .C1(n_0_2447), .C2(n_0_2354), .ZN(n_0_101_2));
   INV_X1 i_0_101_5 (.A(n_0_101_2), .ZN(n_0_2451));
   AOI222_X1 i_0_101_6 (.A1(n_0_2448), .A2(n_0_2418), .B1(n_0_2449), .B2(
      n_0_2386), .C1(n_0_2447), .C2(n_0_2355), .ZN(n_0_101_3));
   INV_X1 i_0_101_7 (.A(n_0_101_3), .ZN(n_0_2452));
   AOI222_X1 i_0_101_8 (.A1(n_0_2448), .A2(n_0_2419), .B1(n_0_2449), .B2(
      n_0_2387), .C1(n_0_2447), .C2(n_0_2356), .ZN(n_0_101_4));
   INV_X1 i_0_101_9 (.A(n_0_101_4), .ZN(n_0_2453));
   AOI222_X1 i_0_101_10 (.A1(n_0_2448), .A2(n_0_2420), .B1(n_0_2449), .B2(
      n_0_2388), .C1(n_0_2447), .C2(n_0_2357), .ZN(n_0_101_5));
   INV_X1 i_0_101_11 (.A(n_0_101_5), .ZN(n_0_2454));
   AOI222_X1 i_0_101_12 (.A1(n_0_2448), .A2(n_0_2421), .B1(n_0_2449), .B2(
      n_0_2389), .C1(n_0_2447), .C2(n_0_2358), .ZN(n_0_101_6));
   INV_X1 i_0_101_13 (.A(n_0_101_6), .ZN(n_0_2455));
   AOI222_X1 i_0_101_14 (.A1(n_0_2448), .A2(n_0_2422), .B1(n_0_2449), .B2(
      n_0_2390), .C1(n_0_2447), .C2(n_0_2359), .ZN(n_0_101_7));
   INV_X1 i_0_101_15 (.A(n_0_101_7), .ZN(n_0_2456));
   AOI222_X1 i_0_101_16 (.A1(n_0_2448), .A2(n_0_2423), .B1(n_0_2449), .B2(
      n_0_2391), .C1(n_0_2447), .C2(n_0_2360), .ZN(n_0_101_8));
   INV_X1 i_0_101_17 (.A(n_0_101_8), .ZN(n_0_2457));
   AOI222_X1 i_0_101_18 (.A1(n_0_2448), .A2(n_0_2424), .B1(n_0_2449), .B2(
      n_0_2392), .C1(n_0_2447), .C2(n_0_2361), .ZN(n_0_101_9));
   INV_X1 i_0_101_19 (.A(n_0_101_9), .ZN(n_0_2458));
   AOI222_X1 i_0_101_20 (.A1(n_0_2448), .A2(n_0_2425), .B1(n_0_2449), .B2(
      n_0_2393), .C1(n_0_2447), .C2(n_0_2362), .ZN(n_0_101_10));
   INV_X1 i_0_101_21 (.A(n_0_101_10), .ZN(n_0_2459));
   AOI222_X1 i_0_101_22 (.A1(n_0_2448), .A2(n_0_2426), .B1(n_0_2449), .B2(
      n_0_2394), .C1(n_0_2447), .C2(n_0_2363), .ZN(n_0_101_11));
   INV_X1 i_0_101_23 (.A(n_0_101_11), .ZN(n_0_2460));
   AOI222_X1 i_0_101_24 (.A1(n_0_2448), .A2(n_0_2427), .B1(n_0_2449), .B2(
      n_0_2395), .C1(n_0_2447), .C2(n_0_2364), .ZN(n_0_101_12));
   INV_X1 i_0_101_25 (.A(n_0_101_12), .ZN(n_0_2461));
   AOI222_X1 i_0_101_26 (.A1(n_0_2448), .A2(n_0_2428), .B1(n_0_2449), .B2(
      n_0_2396), .C1(n_0_2447), .C2(n_0_2365), .ZN(n_0_101_13));
   INV_X1 i_0_101_27 (.A(n_0_101_13), .ZN(n_0_2462));
   AOI222_X1 i_0_101_28 (.A1(n_0_2448), .A2(n_0_2429), .B1(n_0_2449), .B2(
      n_0_2397), .C1(n_0_2447), .C2(n_0_2366), .ZN(n_0_101_14));
   INV_X1 i_0_101_29 (.A(n_0_101_14), .ZN(n_0_2463));
   AOI222_X1 i_0_101_30 (.A1(n_0_2448), .A2(n_0_2430), .B1(n_0_2449), .B2(
      n_0_2398), .C1(n_0_2447), .C2(n_0_2367), .ZN(n_0_101_15));
   INV_X1 i_0_101_31 (.A(n_0_101_15), .ZN(n_0_2464));
   AOI222_X1 i_0_101_32 (.A1(n_0_2448), .A2(n_0_2431), .B1(n_0_2449), .B2(
      n_0_2399), .C1(n_0_2447), .C2(n_0_2368), .ZN(n_0_101_16));
   INV_X1 i_0_101_33 (.A(n_0_101_16), .ZN(n_0_2465));
   AOI222_X1 i_0_101_34 (.A1(n_0_2448), .A2(n_0_2432), .B1(n_0_2449), .B2(
      n_0_2400), .C1(n_0_2447), .C2(n_0_2369), .ZN(n_0_101_17));
   INV_X1 i_0_101_35 (.A(n_0_101_17), .ZN(n_0_2466));
   AOI222_X1 i_0_101_36 (.A1(n_0_2448), .A2(n_0_2433), .B1(n_0_2449), .B2(
      n_0_2401), .C1(n_0_2447), .C2(n_0_2370), .ZN(n_0_101_18));
   INV_X1 i_0_101_37 (.A(n_0_101_18), .ZN(n_0_2467));
   AOI222_X1 i_0_101_38 (.A1(n_0_2448), .A2(n_0_2434), .B1(n_0_2449), .B2(
      n_0_2402), .C1(n_0_2447), .C2(n_0_2371), .ZN(n_0_101_19));
   INV_X1 i_0_101_39 (.A(n_0_101_19), .ZN(n_0_2468));
   AOI222_X1 i_0_101_40 (.A1(n_0_2448), .A2(n_0_2435), .B1(n_0_2449), .B2(
      n_0_2403), .C1(n_0_2447), .C2(n_0_2372), .ZN(n_0_101_20));
   INV_X1 i_0_101_41 (.A(n_0_101_20), .ZN(n_0_2469));
   AOI222_X1 i_0_101_42 (.A1(n_0_2448), .A2(n_0_2436), .B1(n_0_2449), .B2(
      n_0_2404), .C1(n_0_2447), .C2(n_0_2373), .ZN(n_0_101_21));
   INV_X1 i_0_101_43 (.A(n_0_101_21), .ZN(n_0_2470));
   AOI222_X1 i_0_101_44 (.A1(n_0_2448), .A2(n_0_2437), .B1(n_0_2449), .B2(
      n_0_2405), .C1(n_0_2447), .C2(n_0_2374), .ZN(n_0_101_22));
   INV_X1 i_0_101_45 (.A(n_0_101_22), .ZN(n_0_2471));
   AOI222_X1 i_0_101_46 (.A1(n_0_2448), .A2(n_0_2438), .B1(n_0_2449), .B2(
      n_0_2406), .C1(n_0_2447), .C2(n_0_2375), .ZN(n_0_101_23));
   INV_X1 i_0_101_47 (.A(n_0_101_23), .ZN(n_0_2472));
   AOI222_X1 i_0_101_48 (.A1(n_0_2448), .A2(n_0_2439), .B1(n_0_2449), .B2(
      n_0_2407), .C1(n_0_2447), .C2(n_0_2376), .ZN(n_0_101_24));
   INV_X1 i_0_101_49 (.A(n_0_101_24), .ZN(n_0_2473));
   AOI222_X1 i_0_101_50 (.A1(n_0_2448), .A2(n_0_2440), .B1(n_0_2449), .B2(
      n_0_2408), .C1(n_0_2447), .C2(n_0_2377), .ZN(n_0_101_25));
   INV_X1 i_0_101_51 (.A(n_0_101_25), .ZN(n_0_2474));
   AOI222_X1 i_0_101_52 (.A1(n_0_2448), .A2(n_0_2441), .B1(n_0_2449), .B2(
      n_0_2409), .C1(n_0_2447), .C2(n_0_2378), .ZN(n_0_101_26));
   INV_X1 i_0_101_53 (.A(n_0_101_26), .ZN(n_0_2475));
   AOI222_X1 i_0_101_54 (.A1(n_0_2448), .A2(n_0_2442), .B1(n_0_2449), .B2(
      n_0_2410), .C1(n_0_2447), .C2(n_0_2379), .ZN(n_0_101_27));
   INV_X1 i_0_101_55 (.A(n_0_101_27), .ZN(n_0_2476));
   AOI222_X1 i_0_101_56 (.A1(n_0_2448), .A2(n_0_2443), .B1(n_0_2449), .B2(
      n_0_2411), .C1(n_0_2447), .C2(n_0_2380), .ZN(n_0_101_28));
   INV_X1 i_0_101_57 (.A(n_0_101_28), .ZN(n_0_2477));
   AOI222_X1 i_0_101_58 (.A1(n_0_2448), .A2(n_0_2444), .B1(n_0_2449), .B2(
      n_0_2412), .C1(n_0_2447), .C2(n_0_2381), .ZN(n_0_101_29));
   INV_X1 i_0_101_59 (.A(n_0_101_29), .ZN(n_0_2478));
   AND2_X1 i_0_101_60 (.A1(n_0_2447), .A2(n_0_2382), .ZN(n_0_101_30));
   AOI221_X1 i_0_101_61 (.A(n_0_101_30), .B1(n_0_2448), .B2(n_0_2445), .C1(
      n_0_2449), .C2(n_0_2413), .ZN(n_0_101_31));
   INV_X1 i_0_101_62 (.A(n_0_101_31), .ZN(n_0_2479));
   AOI221_X1 i_0_101_63 (.A(n_0_101_30), .B1(n_0_2448), .B2(n_0_2446), .C1(
      n_0_2449), .C2(n_0_2414), .ZN(n_0_101_32));
   INV_X1 i_0_101_64 (.A(n_0_101_32), .ZN(n_0_2480));
   datapath__0_100 i_0_102 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_51, 
      n_0_2480, n_0_2479, n_0_2478, n_0_2477, n_0_2476, n_0_2475, n_0_2474, 
      n_0_2473, n_0_2472, n_0_2471, n_0_2470, n_0_2469, n_0_2468, n_0_2467, 
      n_0_2466, n_0_2465, n_0_2464, n_0_2463, n_0_2462, n_0_2461, n_0_2460, 
      n_0_2459, n_0_2458, n_0_2457, n_0_2456, n_0_2455, n_0_2454, n_0_2453, 
      n_0_2452, n_0_2451, n_0_2450}), .p_2({n_0_2512, n_0_2511, n_0_2510, 
      n_0_2509, n_0_2508, n_0_2507, n_0_2506, n_0_2505, n_0_2504, n_0_2503, 
      n_0_2502, n_0_2501, n_0_2500, n_0_2499, n_0_2498, n_0_2497, n_0_2496, 
      n_0_2495, n_0_2494, n_0_2493, n_0_2492, n_0_2491, n_0_2490, n_0_2489, 
      n_0_2488, n_0_2487, n_0_2486, n_0_2485, n_0_2484, n_0_2483, n_0_2482, 
      n_0_2481}));
   datapath__0_101 i_0_103 (.multiplicand2(multiplicand2), .p_0({uc_52, n_0_2480, 
      n_0_2479, n_0_2478, n_0_2477, n_0_2476, n_0_2475, n_0_2474, n_0_2473, 
      n_0_2472, n_0_2471, n_0_2470, n_0_2469, n_0_2468, n_0_2467, n_0_2466, 
      n_0_2465, n_0_2464, n_0_2463, n_0_2462, n_0_2461, n_0_2460, n_0_2459, 
      n_0_2458, n_0_2457, n_0_2456, n_0_2455, n_0_2454, n_0_2453, n_0_2452, 
      n_0_2451, n_0_2450}), .p_1({n_0_2544, n_0_2543, n_0_2542, n_0_2541, 
      n_0_2540, n_0_2539, n_0_2538, n_0_2537, n_0_2536, n_0_2535, n_0_2534, 
      n_0_2533, n_0_2532, n_0_2531, n_0_2530, n_0_2529, n_0_2528, n_0_2527, 
      n_0_2526, n_0_2525, n_0_2524, n_0_2523, n_0_2522, n_0_2521, n_0_2520, 
      n_0_2519, n_0_2518, n_0_2517, n_0_2516, n_0_2515, n_0_2514, n_0_2513}));
   INV_X1 i_0_104_0 (.A(multiplier2[26]), .ZN(n_0_104_0));
   AND2_X1 i_0_104_1 (.A1(n_0_104_0), .A2(multiplier2[25]), .ZN(n_0_2546));
   NOR2_X1 i_0_104_2 (.A1(n_0_104_0), .A2(multiplier2[25]), .ZN(n_0_2547));
   NOR2_X1 i_0_104_3 (.A1(n_0_2546), .A2(n_0_2547), .ZN(n_0_2545));
   AOI222_X1 i_0_105_0 (.A1(n_0_2513), .A2(n_0_2546), .B1(n_0_2481), .B2(
      n_0_2547), .C1(n_0_2450), .C2(n_0_2545), .ZN(n_0_105_0));
   INV_X1 i_0_105_1 (.A(n_0_105_0), .ZN(product[26]));
   AOI222_X1 i_0_105_2 (.A1(n_0_2546), .A2(n_0_2514), .B1(n_0_2547), .B2(
      n_0_2482), .C1(n_0_2545), .C2(n_0_2451), .ZN(n_0_105_1));
   INV_X1 i_0_105_3 (.A(n_0_105_1), .ZN(n_0_2548));
   AOI222_X1 i_0_105_4 (.A1(n_0_2546), .A2(n_0_2515), .B1(n_0_2547), .B2(
      n_0_2483), .C1(n_0_2545), .C2(n_0_2452), .ZN(n_0_105_2));
   INV_X1 i_0_105_5 (.A(n_0_105_2), .ZN(n_0_2549));
   AOI222_X1 i_0_105_6 (.A1(n_0_2546), .A2(n_0_2516), .B1(n_0_2547), .B2(
      n_0_2484), .C1(n_0_2545), .C2(n_0_2453), .ZN(n_0_105_3));
   INV_X1 i_0_105_7 (.A(n_0_105_3), .ZN(n_0_2550));
   AOI222_X1 i_0_105_8 (.A1(n_0_2546), .A2(n_0_2517), .B1(n_0_2547), .B2(
      n_0_2485), .C1(n_0_2545), .C2(n_0_2454), .ZN(n_0_105_4));
   INV_X1 i_0_105_9 (.A(n_0_105_4), .ZN(n_0_2551));
   AOI222_X1 i_0_105_10 (.A1(n_0_2546), .A2(n_0_2518), .B1(n_0_2547), .B2(
      n_0_2486), .C1(n_0_2545), .C2(n_0_2455), .ZN(n_0_105_5));
   INV_X1 i_0_105_11 (.A(n_0_105_5), .ZN(n_0_2552));
   AOI222_X1 i_0_105_12 (.A1(n_0_2546), .A2(n_0_2519), .B1(n_0_2547), .B2(
      n_0_2487), .C1(n_0_2545), .C2(n_0_2456), .ZN(n_0_105_6));
   INV_X1 i_0_105_13 (.A(n_0_105_6), .ZN(n_0_2553));
   AOI222_X1 i_0_105_14 (.A1(n_0_2546), .A2(n_0_2520), .B1(n_0_2547), .B2(
      n_0_2488), .C1(n_0_2545), .C2(n_0_2457), .ZN(n_0_105_7));
   INV_X1 i_0_105_15 (.A(n_0_105_7), .ZN(n_0_2554));
   AOI222_X1 i_0_105_16 (.A1(n_0_2546), .A2(n_0_2521), .B1(n_0_2547), .B2(
      n_0_2489), .C1(n_0_2545), .C2(n_0_2458), .ZN(n_0_105_8));
   INV_X1 i_0_105_17 (.A(n_0_105_8), .ZN(n_0_2555));
   AOI222_X1 i_0_105_18 (.A1(n_0_2546), .A2(n_0_2522), .B1(n_0_2547), .B2(
      n_0_2490), .C1(n_0_2545), .C2(n_0_2459), .ZN(n_0_105_9));
   INV_X1 i_0_105_19 (.A(n_0_105_9), .ZN(n_0_2556));
   AOI222_X1 i_0_105_20 (.A1(n_0_2546), .A2(n_0_2523), .B1(n_0_2547), .B2(
      n_0_2491), .C1(n_0_2545), .C2(n_0_2460), .ZN(n_0_105_10));
   INV_X1 i_0_105_21 (.A(n_0_105_10), .ZN(n_0_2557));
   AOI222_X1 i_0_105_22 (.A1(n_0_2546), .A2(n_0_2524), .B1(n_0_2547), .B2(
      n_0_2492), .C1(n_0_2545), .C2(n_0_2461), .ZN(n_0_105_11));
   INV_X1 i_0_105_23 (.A(n_0_105_11), .ZN(n_0_2558));
   AOI222_X1 i_0_105_24 (.A1(n_0_2546), .A2(n_0_2525), .B1(n_0_2547), .B2(
      n_0_2493), .C1(n_0_2545), .C2(n_0_2462), .ZN(n_0_105_12));
   INV_X1 i_0_105_25 (.A(n_0_105_12), .ZN(n_0_2559));
   AOI222_X1 i_0_105_26 (.A1(n_0_2546), .A2(n_0_2526), .B1(n_0_2547), .B2(
      n_0_2494), .C1(n_0_2545), .C2(n_0_2463), .ZN(n_0_105_13));
   INV_X1 i_0_105_27 (.A(n_0_105_13), .ZN(n_0_2560));
   AOI222_X1 i_0_105_28 (.A1(n_0_2546), .A2(n_0_2527), .B1(n_0_2547), .B2(
      n_0_2495), .C1(n_0_2545), .C2(n_0_2464), .ZN(n_0_105_14));
   INV_X1 i_0_105_29 (.A(n_0_105_14), .ZN(n_0_2561));
   AOI222_X1 i_0_105_30 (.A1(n_0_2546), .A2(n_0_2528), .B1(n_0_2547), .B2(
      n_0_2496), .C1(n_0_2545), .C2(n_0_2465), .ZN(n_0_105_15));
   INV_X1 i_0_105_31 (.A(n_0_105_15), .ZN(n_0_2562));
   AOI222_X1 i_0_105_32 (.A1(n_0_2546), .A2(n_0_2529), .B1(n_0_2547), .B2(
      n_0_2497), .C1(n_0_2545), .C2(n_0_2466), .ZN(n_0_105_16));
   INV_X1 i_0_105_33 (.A(n_0_105_16), .ZN(n_0_2563));
   AOI222_X1 i_0_105_34 (.A1(n_0_2546), .A2(n_0_2530), .B1(n_0_2547), .B2(
      n_0_2498), .C1(n_0_2545), .C2(n_0_2467), .ZN(n_0_105_17));
   INV_X1 i_0_105_35 (.A(n_0_105_17), .ZN(n_0_2564));
   AOI222_X1 i_0_105_36 (.A1(n_0_2546), .A2(n_0_2531), .B1(n_0_2547), .B2(
      n_0_2499), .C1(n_0_2545), .C2(n_0_2468), .ZN(n_0_105_18));
   INV_X1 i_0_105_37 (.A(n_0_105_18), .ZN(n_0_2565));
   AOI222_X1 i_0_105_38 (.A1(n_0_2546), .A2(n_0_2532), .B1(n_0_2547), .B2(
      n_0_2500), .C1(n_0_2545), .C2(n_0_2469), .ZN(n_0_105_19));
   INV_X1 i_0_105_39 (.A(n_0_105_19), .ZN(n_0_2566));
   AOI222_X1 i_0_105_40 (.A1(n_0_2546), .A2(n_0_2533), .B1(n_0_2547), .B2(
      n_0_2501), .C1(n_0_2545), .C2(n_0_2470), .ZN(n_0_105_20));
   INV_X1 i_0_105_41 (.A(n_0_105_20), .ZN(n_0_2567));
   AOI222_X1 i_0_105_42 (.A1(n_0_2546), .A2(n_0_2534), .B1(n_0_2547), .B2(
      n_0_2502), .C1(n_0_2545), .C2(n_0_2471), .ZN(n_0_105_21));
   INV_X1 i_0_105_43 (.A(n_0_105_21), .ZN(n_0_2568));
   AOI222_X1 i_0_105_44 (.A1(n_0_2546), .A2(n_0_2535), .B1(n_0_2547), .B2(
      n_0_2503), .C1(n_0_2545), .C2(n_0_2472), .ZN(n_0_105_22));
   INV_X1 i_0_105_45 (.A(n_0_105_22), .ZN(n_0_2569));
   AOI222_X1 i_0_105_46 (.A1(n_0_2546), .A2(n_0_2536), .B1(n_0_2547), .B2(
      n_0_2504), .C1(n_0_2545), .C2(n_0_2473), .ZN(n_0_105_23));
   INV_X1 i_0_105_47 (.A(n_0_105_23), .ZN(n_0_2570));
   AOI222_X1 i_0_105_48 (.A1(n_0_2546), .A2(n_0_2537), .B1(n_0_2547), .B2(
      n_0_2505), .C1(n_0_2545), .C2(n_0_2474), .ZN(n_0_105_24));
   INV_X1 i_0_105_49 (.A(n_0_105_24), .ZN(n_0_2571));
   AOI222_X1 i_0_105_50 (.A1(n_0_2546), .A2(n_0_2538), .B1(n_0_2547), .B2(
      n_0_2506), .C1(n_0_2545), .C2(n_0_2475), .ZN(n_0_105_25));
   INV_X1 i_0_105_51 (.A(n_0_105_25), .ZN(n_0_2572));
   AOI222_X1 i_0_105_52 (.A1(n_0_2546), .A2(n_0_2539), .B1(n_0_2547), .B2(
      n_0_2507), .C1(n_0_2545), .C2(n_0_2476), .ZN(n_0_105_26));
   INV_X1 i_0_105_53 (.A(n_0_105_26), .ZN(n_0_2573));
   AOI222_X1 i_0_105_54 (.A1(n_0_2546), .A2(n_0_2540), .B1(n_0_2547), .B2(
      n_0_2508), .C1(n_0_2545), .C2(n_0_2477), .ZN(n_0_105_27));
   INV_X1 i_0_105_55 (.A(n_0_105_27), .ZN(n_0_2574));
   AOI222_X1 i_0_105_56 (.A1(n_0_2546), .A2(n_0_2541), .B1(n_0_2547), .B2(
      n_0_2509), .C1(n_0_2545), .C2(n_0_2478), .ZN(n_0_105_28));
   INV_X1 i_0_105_57 (.A(n_0_105_28), .ZN(n_0_2575));
   AOI222_X1 i_0_105_58 (.A1(n_0_2546), .A2(n_0_2542), .B1(n_0_2547), .B2(
      n_0_2510), .C1(n_0_2545), .C2(n_0_2479), .ZN(n_0_105_29));
   INV_X1 i_0_105_59 (.A(n_0_105_29), .ZN(n_0_2576));
   AND2_X1 i_0_105_60 (.A1(n_0_2545), .A2(n_0_2480), .ZN(n_0_105_30));
   AOI221_X1 i_0_105_61 (.A(n_0_105_30), .B1(n_0_2546), .B2(n_0_2543), .C1(
      n_0_2547), .C2(n_0_2511), .ZN(n_0_105_31));
   INV_X1 i_0_105_62 (.A(n_0_105_31), .ZN(n_0_2577));
   AOI221_X1 i_0_105_63 (.A(n_0_105_30), .B1(n_0_2546), .B2(n_0_2544), .C1(
      n_0_2547), .C2(n_0_2512), .ZN(n_0_105_32));
   INV_X1 i_0_105_64 (.A(n_0_105_32), .ZN(n_0_2578));
   datapath__0_104 i_0_106 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_53, 
      n_0_2578, n_0_2577, n_0_2576, n_0_2575, n_0_2574, n_0_2573, n_0_2572, 
      n_0_2571, n_0_2570, n_0_2569, n_0_2568, n_0_2567, n_0_2566, n_0_2565, 
      n_0_2564, n_0_2563, n_0_2562, n_0_2561, n_0_2560, n_0_2559, n_0_2558, 
      n_0_2557, n_0_2556, n_0_2555, n_0_2554, n_0_2553, n_0_2552, n_0_2551, 
      n_0_2550, n_0_2549, n_0_2548}), .p_2({n_0_2610, n_0_2609, n_0_2608, 
      n_0_2607, n_0_2606, n_0_2605, n_0_2604, n_0_2603, n_0_2602, n_0_2601, 
      n_0_2600, n_0_2599, n_0_2598, n_0_2597, n_0_2596, n_0_2595, n_0_2594, 
      n_0_2593, n_0_2592, n_0_2591, n_0_2590, n_0_2589, n_0_2588, n_0_2587, 
      n_0_2586, n_0_2585, n_0_2584, n_0_2583, n_0_2582, n_0_2581, n_0_2580, 
      n_0_2579}));
   datapath__0_105 i_0_107 (.multiplicand2(multiplicand2), .p_0({uc_54, n_0_2578, 
      n_0_2577, n_0_2576, n_0_2575, n_0_2574, n_0_2573, n_0_2572, n_0_2571, 
      n_0_2570, n_0_2569, n_0_2568, n_0_2567, n_0_2566, n_0_2565, n_0_2564, 
      n_0_2563, n_0_2562, n_0_2561, n_0_2560, n_0_2559, n_0_2558, n_0_2557, 
      n_0_2556, n_0_2555, n_0_2554, n_0_2553, n_0_2552, n_0_2551, n_0_2550, 
      n_0_2549, n_0_2548}), .p_1({n_0_2642, n_0_2641, n_0_2640, n_0_2639, 
      n_0_2638, n_0_2637, n_0_2636, n_0_2635, n_0_2634, n_0_2633, n_0_2632, 
      n_0_2631, n_0_2630, n_0_2629, n_0_2628, n_0_2627, n_0_2626, n_0_2625, 
      n_0_2624, n_0_2623, n_0_2622, n_0_2621, n_0_2620, n_0_2619, n_0_2618, 
      n_0_2617, n_0_2616, n_0_2615, n_0_2614, n_0_2613, n_0_2612, n_0_2611}));
   INV_X1 i_0_108_0 (.A(multiplier2[27]), .ZN(n_0_108_0));
   AND2_X1 i_0_108_1 (.A1(n_0_108_0), .A2(multiplier2[26]), .ZN(n_0_2644));
   NOR2_X1 i_0_108_2 (.A1(n_0_108_0), .A2(multiplier2[26]), .ZN(n_0_2645));
   NOR2_X1 i_0_108_3 (.A1(n_0_2644), .A2(n_0_2645), .ZN(n_0_2643));
   AOI222_X1 i_0_109_0 (.A1(n_0_2611), .A2(n_0_2644), .B1(n_0_2579), .B2(
      n_0_2645), .C1(n_0_2548), .C2(n_0_2643), .ZN(n_0_109_0));
   INV_X1 i_0_109_1 (.A(n_0_109_0), .ZN(product[27]));
   AOI222_X1 i_0_109_2 (.A1(n_0_2644), .A2(n_0_2612), .B1(n_0_2645), .B2(
      n_0_2580), .C1(n_0_2643), .C2(n_0_2549), .ZN(n_0_109_1));
   INV_X1 i_0_109_3 (.A(n_0_109_1), .ZN(n_0_2646));
   AOI222_X1 i_0_109_4 (.A1(n_0_2644), .A2(n_0_2613), .B1(n_0_2645), .B2(
      n_0_2581), .C1(n_0_2643), .C2(n_0_2550), .ZN(n_0_109_2));
   INV_X1 i_0_109_5 (.A(n_0_109_2), .ZN(n_0_2647));
   AOI222_X1 i_0_109_6 (.A1(n_0_2644), .A2(n_0_2614), .B1(n_0_2645), .B2(
      n_0_2582), .C1(n_0_2643), .C2(n_0_2551), .ZN(n_0_109_3));
   INV_X1 i_0_109_7 (.A(n_0_109_3), .ZN(n_0_2648));
   AOI222_X1 i_0_109_8 (.A1(n_0_2644), .A2(n_0_2615), .B1(n_0_2645), .B2(
      n_0_2583), .C1(n_0_2643), .C2(n_0_2552), .ZN(n_0_109_4));
   INV_X1 i_0_109_9 (.A(n_0_109_4), .ZN(n_0_2649));
   AOI222_X1 i_0_109_10 (.A1(n_0_2644), .A2(n_0_2616), .B1(n_0_2645), .B2(
      n_0_2584), .C1(n_0_2643), .C2(n_0_2553), .ZN(n_0_109_5));
   INV_X1 i_0_109_11 (.A(n_0_109_5), .ZN(n_0_2650));
   AOI222_X1 i_0_109_12 (.A1(n_0_2644), .A2(n_0_2617), .B1(n_0_2645), .B2(
      n_0_2585), .C1(n_0_2643), .C2(n_0_2554), .ZN(n_0_109_6));
   INV_X1 i_0_109_13 (.A(n_0_109_6), .ZN(n_0_2651));
   AOI222_X1 i_0_109_14 (.A1(n_0_2644), .A2(n_0_2618), .B1(n_0_2645), .B2(
      n_0_2586), .C1(n_0_2643), .C2(n_0_2555), .ZN(n_0_109_7));
   INV_X1 i_0_109_15 (.A(n_0_109_7), .ZN(n_0_2652));
   AOI222_X1 i_0_109_16 (.A1(n_0_2644), .A2(n_0_2619), .B1(n_0_2645), .B2(
      n_0_2587), .C1(n_0_2643), .C2(n_0_2556), .ZN(n_0_109_8));
   INV_X1 i_0_109_17 (.A(n_0_109_8), .ZN(n_0_2653));
   AOI222_X1 i_0_109_18 (.A1(n_0_2644), .A2(n_0_2620), .B1(n_0_2645), .B2(
      n_0_2588), .C1(n_0_2643), .C2(n_0_2557), .ZN(n_0_109_9));
   INV_X1 i_0_109_19 (.A(n_0_109_9), .ZN(n_0_2654));
   AOI222_X1 i_0_109_20 (.A1(n_0_2644), .A2(n_0_2621), .B1(n_0_2645), .B2(
      n_0_2589), .C1(n_0_2643), .C2(n_0_2558), .ZN(n_0_109_10));
   INV_X1 i_0_109_21 (.A(n_0_109_10), .ZN(n_0_2655));
   AOI222_X1 i_0_109_22 (.A1(n_0_2644), .A2(n_0_2622), .B1(n_0_2645), .B2(
      n_0_2590), .C1(n_0_2643), .C2(n_0_2559), .ZN(n_0_109_11));
   INV_X1 i_0_109_23 (.A(n_0_109_11), .ZN(n_0_2656));
   AOI222_X1 i_0_109_24 (.A1(n_0_2644), .A2(n_0_2623), .B1(n_0_2645), .B2(
      n_0_2591), .C1(n_0_2643), .C2(n_0_2560), .ZN(n_0_109_12));
   INV_X1 i_0_109_25 (.A(n_0_109_12), .ZN(n_0_2657));
   AOI222_X1 i_0_109_26 (.A1(n_0_2644), .A2(n_0_2624), .B1(n_0_2645), .B2(
      n_0_2592), .C1(n_0_2643), .C2(n_0_2561), .ZN(n_0_109_13));
   INV_X1 i_0_109_27 (.A(n_0_109_13), .ZN(n_0_2658));
   AOI222_X1 i_0_109_28 (.A1(n_0_2644), .A2(n_0_2625), .B1(n_0_2645), .B2(
      n_0_2593), .C1(n_0_2643), .C2(n_0_2562), .ZN(n_0_109_14));
   INV_X1 i_0_109_29 (.A(n_0_109_14), .ZN(n_0_2659));
   AOI222_X1 i_0_109_30 (.A1(n_0_2644), .A2(n_0_2626), .B1(n_0_2645), .B2(
      n_0_2594), .C1(n_0_2643), .C2(n_0_2563), .ZN(n_0_109_15));
   INV_X1 i_0_109_31 (.A(n_0_109_15), .ZN(n_0_2660));
   AOI222_X1 i_0_109_32 (.A1(n_0_2644), .A2(n_0_2627), .B1(n_0_2645), .B2(
      n_0_2595), .C1(n_0_2643), .C2(n_0_2564), .ZN(n_0_109_16));
   INV_X1 i_0_109_33 (.A(n_0_109_16), .ZN(n_0_2661));
   AOI222_X1 i_0_109_34 (.A1(n_0_2644), .A2(n_0_2628), .B1(n_0_2645), .B2(
      n_0_2596), .C1(n_0_2643), .C2(n_0_2565), .ZN(n_0_109_17));
   INV_X1 i_0_109_35 (.A(n_0_109_17), .ZN(n_0_2662));
   AOI222_X1 i_0_109_36 (.A1(n_0_2644), .A2(n_0_2629), .B1(n_0_2645), .B2(
      n_0_2597), .C1(n_0_2643), .C2(n_0_2566), .ZN(n_0_109_18));
   INV_X1 i_0_109_37 (.A(n_0_109_18), .ZN(n_0_2663));
   AOI222_X1 i_0_109_38 (.A1(n_0_2644), .A2(n_0_2630), .B1(n_0_2645), .B2(
      n_0_2598), .C1(n_0_2643), .C2(n_0_2567), .ZN(n_0_109_19));
   INV_X1 i_0_109_39 (.A(n_0_109_19), .ZN(n_0_2664));
   AOI222_X1 i_0_109_40 (.A1(n_0_2644), .A2(n_0_2631), .B1(n_0_2645), .B2(
      n_0_2599), .C1(n_0_2643), .C2(n_0_2568), .ZN(n_0_109_20));
   INV_X1 i_0_109_41 (.A(n_0_109_20), .ZN(n_0_2665));
   AOI222_X1 i_0_109_42 (.A1(n_0_2644), .A2(n_0_2632), .B1(n_0_2645), .B2(
      n_0_2600), .C1(n_0_2643), .C2(n_0_2569), .ZN(n_0_109_21));
   INV_X1 i_0_109_43 (.A(n_0_109_21), .ZN(n_0_2666));
   AOI222_X1 i_0_109_44 (.A1(n_0_2644), .A2(n_0_2633), .B1(n_0_2645), .B2(
      n_0_2601), .C1(n_0_2643), .C2(n_0_2570), .ZN(n_0_109_22));
   INV_X1 i_0_109_45 (.A(n_0_109_22), .ZN(n_0_2667));
   AOI222_X1 i_0_109_46 (.A1(n_0_2644), .A2(n_0_2634), .B1(n_0_2645), .B2(
      n_0_2602), .C1(n_0_2643), .C2(n_0_2571), .ZN(n_0_109_23));
   INV_X1 i_0_109_47 (.A(n_0_109_23), .ZN(n_0_2668));
   AOI222_X1 i_0_109_48 (.A1(n_0_2644), .A2(n_0_2635), .B1(n_0_2645), .B2(
      n_0_2603), .C1(n_0_2643), .C2(n_0_2572), .ZN(n_0_109_24));
   INV_X1 i_0_109_49 (.A(n_0_109_24), .ZN(n_0_2669));
   AOI222_X1 i_0_109_50 (.A1(n_0_2644), .A2(n_0_2636), .B1(n_0_2645), .B2(
      n_0_2604), .C1(n_0_2643), .C2(n_0_2573), .ZN(n_0_109_25));
   INV_X1 i_0_109_51 (.A(n_0_109_25), .ZN(n_0_2670));
   AOI222_X1 i_0_109_52 (.A1(n_0_2644), .A2(n_0_2637), .B1(n_0_2645), .B2(
      n_0_2605), .C1(n_0_2643), .C2(n_0_2574), .ZN(n_0_109_26));
   INV_X1 i_0_109_53 (.A(n_0_109_26), .ZN(n_0_2671));
   AOI222_X1 i_0_109_54 (.A1(n_0_2644), .A2(n_0_2638), .B1(n_0_2645), .B2(
      n_0_2606), .C1(n_0_2643), .C2(n_0_2575), .ZN(n_0_109_27));
   INV_X1 i_0_109_55 (.A(n_0_109_27), .ZN(n_0_2672));
   AOI222_X1 i_0_109_56 (.A1(n_0_2644), .A2(n_0_2639), .B1(n_0_2645), .B2(
      n_0_2607), .C1(n_0_2643), .C2(n_0_2576), .ZN(n_0_109_28));
   INV_X1 i_0_109_57 (.A(n_0_109_28), .ZN(n_0_2673));
   AOI222_X1 i_0_109_58 (.A1(n_0_2644), .A2(n_0_2640), .B1(n_0_2645), .B2(
      n_0_2608), .C1(n_0_2643), .C2(n_0_2577), .ZN(n_0_109_29));
   INV_X1 i_0_109_59 (.A(n_0_109_29), .ZN(n_0_2674));
   AND2_X1 i_0_109_60 (.A1(n_0_2643), .A2(n_0_2578), .ZN(n_0_109_30));
   AOI221_X1 i_0_109_61 (.A(n_0_109_30), .B1(n_0_2644), .B2(n_0_2641), .C1(
      n_0_2645), .C2(n_0_2609), .ZN(n_0_109_31));
   INV_X1 i_0_109_62 (.A(n_0_109_31), .ZN(n_0_2675));
   AOI221_X1 i_0_109_63 (.A(n_0_109_30), .B1(n_0_2644), .B2(n_0_2642), .C1(
      n_0_2645), .C2(n_0_2610), .ZN(n_0_109_32));
   INV_X1 i_0_109_64 (.A(n_0_109_32), .ZN(n_0_2676));
   datapath__0_108 i_0_110 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_55, 
      n_0_2676, n_0_2675, n_0_2674, n_0_2673, n_0_2672, n_0_2671, n_0_2670, 
      n_0_2669, n_0_2668, n_0_2667, n_0_2666, n_0_2665, n_0_2664, n_0_2663, 
      n_0_2662, n_0_2661, n_0_2660, n_0_2659, n_0_2658, n_0_2657, n_0_2656, 
      n_0_2655, n_0_2654, n_0_2653, n_0_2652, n_0_2651, n_0_2650, n_0_2649, 
      n_0_2648, n_0_2647, n_0_2646}), .p_2({n_0_2708, n_0_2707, n_0_2706, 
      n_0_2705, n_0_2704, n_0_2703, n_0_2702, n_0_2701, n_0_2700, n_0_2699, 
      n_0_2698, n_0_2697, n_0_2696, n_0_2695, n_0_2694, n_0_2693, n_0_2692, 
      n_0_2691, n_0_2690, n_0_2689, n_0_2688, n_0_2687, n_0_2686, n_0_2685, 
      n_0_2684, n_0_2683, n_0_2682, n_0_2681, n_0_2680, n_0_2679, n_0_2678, 
      n_0_2677}));
   datapath__0_109 i_0_111 (.multiplicand2(multiplicand2), .p_0({uc_56, n_0_2676, 
      n_0_2675, n_0_2674, n_0_2673, n_0_2672, n_0_2671, n_0_2670, n_0_2669, 
      n_0_2668, n_0_2667, n_0_2666, n_0_2665, n_0_2664, n_0_2663, n_0_2662, 
      n_0_2661, n_0_2660, n_0_2659, n_0_2658, n_0_2657, n_0_2656, n_0_2655, 
      n_0_2654, n_0_2653, n_0_2652, n_0_2651, n_0_2650, n_0_2649, n_0_2648, 
      n_0_2647, n_0_2646}), .p_1({n_0_2740, n_0_2739, n_0_2738, n_0_2737, 
      n_0_2736, n_0_2735, n_0_2734, n_0_2733, n_0_2732, n_0_2731, n_0_2730, 
      n_0_2729, n_0_2728, n_0_2727, n_0_2726, n_0_2725, n_0_2724, n_0_2723, 
      n_0_2722, n_0_2721, n_0_2720, n_0_2719, n_0_2718, n_0_2717, n_0_2716, 
      n_0_2715, n_0_2714, n_0_2713, n_0_2712, n_0_2711, n_0_2710, n_0_2709}));
   INV_X1 i_0_112_0 (.A(multiplier2[28]), .ZN(n_0_112_0));
   AND2_X1 i_0_112_1 (.A1(n_0_112_0), .A2(multiplier2[27]), .ZN(n_0_2742));
   NOR2_X1 i_0_112_2 (.A1(n_0_112_0), .A2(multiplier2[27]), .ZN(n_0_2743));
   NOR2_X1 i_0_112_3 (.A1(n_0_2742), .A2(n_0_2743), .ZN(n_0_2741));
   AOI222_X1 i_0_113_0 (.A1(n_0_2709), .A2(n_0_2742), .B1(n_0_2677), .B2(
      n_0_2743), .C1(n_0_2646), .C2(n_0_2741), .ZN(n_0_113_0));
   INV_X1 i_0_113_1 (.A(n_0_113_0), .ZN(product[28]));
   AOI222_X1 i_0_113_2 (.A1(n_0_2742), .A2(n_0_2710), .B1(n_0_2743), .B2(
      n_0_2678), .C1(n_0_2741), .C2(n_0_2647), .ZN(n_0_113_1));
   INV_X1 i_0_113_3 (.A(n_0_113_1), .ZN(n_0_2744));
   AOI222_X1 i_0_113_4 (.A1(n_0_2742), .A2(n_0_2711), .B1(n_0_2743), .B2(
      n_0_2679), .C1(n_0_2741), .C2(n_0_2648), .ZN(n_0_113_2));
   INV_X1 i_0_113_5 (.A(n_0_113_2), .ZN(n_0_2745));
   AOI222_X1 i_0_113_6 (.A1(n_0_2742), .A2(n_0_2712), .B1(n_0_2743), .B2(
      n_0_2680), .C1(n_0_2741), .C2(n_0_2649), .ZN(n_0_113_3));
   INV_X1 i_0_113_7 (.A(n_0_113_3), .ZN(n_0_2746));
   AOI222_X1 i_0_113_8 (.A1(n_0_2742), .A2(n_0_2713), .B1(n_0_2743), .B2(
      n_0_2681), .C1(n_0_2741), .C2(n_0_2650), .ZN(n_0_113_4));
   INV_X1 i_0_113_9 (.A(n_0_113_4), .ZN(n_0_2747));
   AOI222_X1 i_0_113_10 (.A1(n_0_2742), .A2(n_0_2714), .B1(n_0_2743), .B2(
      n_0_2682), .C1(n_0_2741), .C2(n_0_2651), .ZN(n_0_113_5));
   INV_X1 i_0_113_11 (.A(n_0_113_5), .ZN(n_0_2748));
   AOI222_X1 i_0_113_12 (.A1(n_0_2742), .A2(n_0_2715), .B1(n_0_2743), .B2(
      n_0_2683), .C1(n_0_2741), .C2(n_0_2652), .ZN(n_0_113_6));
   INV_X1 i_0_113_13 (.A(n_0_113_6), .ZN(n_0_2749));
   AOI222_X1 i_0_113_14 (.A1(n_0_2742), .A2(n_0_2716), .B1(n_0_2743), .B2(
      n_0_2684), .C1(n_0_2741), .C2(n_0_2653), .ZN(n_0_113_7));
   INV_X1 i_0_113_15 (.A(n_0_113_7), .ZN(n_0_2750));
   AOI222_X1 i_0_113_16 (.A1(n_0_2742), .A2(n_0_2717), .B1(n_0_2743), .B2(
      n_0_2685), .C1(n_0_2741), .C2(n_0_2654), .ZN(n_0_113_8));
   INV_X1 i_0_113_17 (.A(n_0_113_8), .ZN(n_0_2751));
   AOI222_X1 i_0_113_18 (.A1(n_0_2742), .A2(n_0_2718), .B1(n_0_2743), .B2(
      n_0_2686), .C1(n_0_2741), .C2(n_0_2655), .ZN(n_0_113_9));
   INV_X1 i_0_113_19 (.A(n_0_113_9), .ZN(n_0_2752));
   AOI222_X1 i_0_113_20 (.A1(n_0_2742), .A2(n_0_2719), .B1(n_0_2743), .B2(
      n_0_2687), .C1(n_0_2741), .C2(n_0_2656), .ZN(n_0_113_10));
   INV_X1 i_0_113_21 (.A(n_0_113_10), .ZN(n_0_2753));
   AOI222_X1 i_0_113_22 (.A1(n_0_2742), .A2(n_0_2720), .B1(n_0_2743), .B2(
      n_0_2688), .C1(n_0_2741), .C2(n_0_2657), .ZN(n_0_113_11));
   INV_X1 i_0_113_23 (.A(n_0_113_11), .ZN(n_0_2754));
   AOI222_X1 i_0_113_24 (.A1(n_0_2742), .A2(n_0_2721), .B1(n_0_2743), .B2(
      n_0_2689), .C1(n_0_2741), .C2(n_0_2658), .ZN(n_0_113_12));
   INV_X1 i_0_113_25 (.A(n_0_113_12), .ZN(n_0_2755));
   AOI222_X1 i_0_113_26 (.A1(n_0_2742), .A2(n_0_2722), .B1(n_0_2743), .B2(
      n_0_2690), .C1(n_0_2741), .C2(n_0_2659), .ZN(n_0_113_13));
   INV_X1 i_0_113_27 (.A(n_0_113_13), .ZN(n_0_2756));
   AOI222_X1 i_0_113_28 (.A1(n_0_2742), .A2(n_0_2723), .B1(n_0_2743), .B2(
      n_0_2691), .C1(n_0_2741), .C2(n_0_2660), .ZN(n_0_113_14));
   INV_X1 i_0_113_29 (.A(n_0_113_14), .ZN(n_0_2757));
   AOI222_X1 i_0_113_30 (.A1(n_0_2742), .A2(n_0_2724), .B1(n_0_2743), .B2(
      n_0_2692), .C1(n_0_2741), .C2(n_0_2661), .ZN(n_0_113_15));
   INV_X1 i_0_113_31 (.A(n_0_113_15), .ZN(n_0_2758));
   AOI222_X1 i_0_113_32 (.A1(n_0_2742), .A2(n_0_2725), .B1(n_0_2743), .B2(
      n_0_2693), .C1(n_0_2741), .C2(n_0_2662), .ZN(n_0_113_16));
   INV_X1 i_0_113_33 (.A(n_0_113_16), .ZN(n_0_2759));
   AOI222_X1 i_0_113_34 (.A1(n_0_2742), .A2(n_0_2726), .B1(n_0_2743), .B2(
      n_0_2694), .C1(n_0_2741), .C2(n_0_2663), .ZN(n_0_113_17));
   INV_X1 i_0_113_35 (.A(n_0_113_17), .ZN(n_0_2760));
   AOI222_X1 i_0_113_36 (.A1(n_0_2742), .A2(n_0_2727), .B1(n_0_2743), .B2(
      n_0_2695), .C1(n_0_2741), .C2(n_0_2664), .ZN(n_0_113_18));
   INV_X1 i_0_113_37 (.A(n_0_113_18), .ZN(n_0_2761));
   AOI222_X1 i_0_113_38 (.A1(n_0_2742), .A2(n_0_2728), .B1(n_0_2743), .B2(
      n_0_2696), .C1(n_0_2741), .C2(n_0_2665), .ZN(n_0_113_19));
   INV_X1 i_0_113_39 (.A(n_0_113_19), .ZN(n_0_2762));
   AOI222_X1 i_0_113_40 (.A1(n_0_2742), .A2(n_0_2729), .B1(n_0_2743), .B2(
      n_0_2697), .C1(n_0_2741), .C2(n_0_2666), .ZN(n_0_113_20));
   INV_X1 i_0_113_41 (.A(n_0_113_20), .ZN(n_0_2763));
   AOI222_X1 i_0_113_42 (.A1(n_0_2742), .A2(n_0_2730), .B1(n_0_2743), .B2(
      n_0_2698), .C1(n_0_2741), .C2(n_0_2667), .ZN(n_0_113_21));
   INV_X1 i_0_113_43 (.A(n_0_113_21), .ZN(n_0_2764));
   AOI222_X1 i_0_113_44 (.A1(n_0_2742), .A2(n_0_2731), .B1(n_0_2743), .B2(
      n_0_2699), .C1(n_0_2741), .C2(n_0_2668), .ZN(n_0_113_22));
   INV_X1 i_0_113_45 (.A(n_0_113_22), .ZN(n_0_2765));
   AOI222_X1 i_0_113_46 (.A1(n_0_2742), .A2(n_0_2732), .B1(n_0_2743), .B2(
      n_0_2700), .C1(n_0_2741), .C2(n_0_2669), .ZN(n_0_113_23));
   INV_X1 i_0_113_47 (.A(n_0_113_23), .ZN(n_0_2766));
   AOI222_X1 i_0_113_48 (.A1(n_0_2742), .A2(n_0_2733), .B1(n_0_2743), .B2(
      n_0_2701), .C1(n_0_2741), .C2(n_0_2670), .ZN(n_0_113_24));
   INV_X1 i_0_113_49 (.A(n_0_113_24), .ZN(n_0_2767));
   AOI222_X1 i_0_113_50 (.A1(n_0_2742), .A2(n_0_2734), .B1(n_0_2743), .B2(
      n_0_2702), .C1(n_0_2741), .C2(n_0_2671), .ZN(n_0_113_25));
   INV_X1 i_0_113_51 (.A(n_0_113_25), .ZN(n_0_2768));
   AOI222_X1 i_0_113_52 (.A1(n_0_2742), .A2(n_0_2735), .B1(n_0_2743), .B2(
      n_0_2703), .C1(n_0_2741), .C2(n_0_2672), .ZN(n_0_113_26));
   INV_X1 i_0_113_53 (.A(n_0_113_26), .ZN(n_0_2769));
   AOI222_X1 i_0_113_54 (.A1(n_0_2742), .A2(n_0_2736), .B1(n_0_2743), .B2(
      n_0_2704), .C1(n_0_2741), .C2(n_0_2673), .ZN(n_0_113_27));
   INV_X1 i_0_113_55 (.A(n_0_113_27), .ZN(n_0_2770));
   AOI222_X1 i_0_113_56 (.A1(n_0_2742), .A2(n_0_2737), .B1(n_0_2743), .B2(
      n_0_2705), .C1(n_0_2741), .C2(n_0_2674), .ZN(n_0_113_28));
   INV_X1 i_0_113_57 (.A(n_0_113_28), .ZN(n_0_2771));
   AOI222_X1 i_0_113_58 (.A1(n_0_2742), .A2(n_0_2738), .B1(n_0_2743), .B2(
      n_0_2706), .C1(n_0_2741), .C2(n_0_2675), .ZN(n_0_113_29));
   INV_X1 i_0_113_59 (.A(n_0_113_29), .ZN(n_0_2772));
   AND2_X1 i_0_113_60 (.A1(n_0_2741), .A2(n_0_2676), .ZN(n_0_113_30));
   AOI221_X1 i_0_113_61 (.A(n_0_113_30), .B1(n_0_2742), .B2(n_0_2739), .C1(
      n_0_2743), .C2(n_0_2707), .ZN(n_0_113_31));
   INV_X1 i_0_113_62 (.A(n_0_113_31), .ZN(n_0_2773));
   AOI221_X1 i_0_113_63 (.A(n_0_113_30), .B1(n_0_2742), .B2(n_0_2740), .C1(
      n_0_2743), .C2(n_0_2708), .ZN(n_0_113_32));
   INV_X1 i_0_113_64 (.A(n_0_113_32), .ZN(n_0_2774));
   datapath__0_112 i_0_114 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_57, 
      n_0_2774, n_0_2773, n_0_2772, n_0_2771, n_0_2770, n_0_2769, n_0_2768, 
      n_0_2767, n_0_2766, n_0_2765, n_0_2764, n_0_2763, n_0_2762, n_0_2761, 
      n_0_2760, n_0_2759, n_0_2758, n_0_2757, n_0_2756, n_0_2755, n_0_2754, 
      n_0_2753, n_0_2752, n_0_2751, n_0_2750, n_0_2749, n_0_2748, n_0_2747, 
      n_0_2746, n_0_2745, n_0_2744}), .p_2({n_0_2806, n_0_2805, n_0_2804, 
      n_0_2803, n_0_2802, n_0_2801, n_0_2800, n_0_2799, n_0_2798, n_0_2797, 
      n_0_2796, n_0_2795, n_0_2794, n_0_2793, n_0_2792, n_0_2791, n_0_2790, 
      n_0_2789, n_0_2788, n_0_2787, n_0_2786, n_0_2785, n_0_2784, n_0_2783, 
      n_0_2782, n_0_2781, n_0_2780, n_0_2779, n_0_2778, n_0_2777, n_0_2776, 
      n_0_2775}));
   datapath__0_113 i_0_115 (.multiplicand2(multiplicand2), .p_0({uc_58, n_0_2774, 
      n_0_2773, n_0_2772, n_0_2771, n_0_2770, n_0_2769, n_0_2768, n_0_2767, 
      n_0_2766, n_0_2765, n_0_2764, n_0_2763, n_0_2762, n_0_2761, n_0_2760, 
      n_0_2759, n_0_2758, n_0_2757, n_0_2756, n_0_2755, n_0_2754, n_0_2753, 
      n_0_2752, n_0_2751, n_0_2750, n_0_2749, n_0_2748, n_0_2747, n_0_2746, 
      n_0_2745, n_0_2744}), .p_1({n_0_2838, n_0_2837, n_0_2836, n_0_2835, 
      n_0_2834, n_0_2833, n_0_2832, n_0_2831, n_0_2830, n_0_2829, n_0_2828, 
      n_0_2827, n_0_2826, n_0_2825, n_0_2824, n_0_2823, n_0_2822, n_0_2821, 
      n_0_2820, n_0_2819, n_0_2818, n_0_2817, n_0_2816, n_0_2815, n_0_2814, 
      n_0_2813, n_0_2812, n_0_2811, n_0_2810, n_0_2809, n_0_2808, n_0_2807}));
   INV_X1 i_0_116_0 (.A(multiplier2[29]), .ZN(n_0_116_0));
   AND2_X1 i_0_116_1 (.A1(n_0_116_0), .A2(multiplier2[28]), .ZN(n_0_2840));
   NOR2_X1 i_0_116_2 (.A1(n_0_116_0), .A2(multiplier2[28]), .ZN(n_0_2841));
   NOR2_X1 i_0_116_3 (.A1(n_0_2840), .A2(n_0_2841), .ZN(n_0_2839));
   AOI222_X1 i_0_117_0 (.A1(n_0_2807), .A2(n_0_2840), .B1(n_0_2775), .B2(
      n_0_2841), .C1(n_0_2744), .C2(n_0_2839), .ZN(n_0_117_0));
   INV_X1 i_0_117_1 (.A(n_0_117_0), .ZN(product[29]));
   AOI222_X1 i_0_117_2 (.A1(n_0_2840), .A2(n_0_2808), .B1(n_0_2841), .B2(
      n_0_2776), .C1(n_0_2839), .C2(n_0_2745), .ZN(n_0_117_1));
   INV_X1 i_0_117_3 (.A(n_0_117_1), .ZN(n_0_2842));
   AOI222_X1 i_0_117_4 (.A1(n_0_2840), .A2(n_0_2809), .B1(n_0_2841), .B2(
      n_0_2777), .C1(n_0_2839), .C2(n_0_2746), .ZN(n_0_117_2));
   INV_X1 i_0_117_5 (.A(n_0_117_2), .ZN(n_0_2843));
   AOI222_X1 i_0_117_6 (.A1(n_0_2840), .A2(n_0_2810), .B1(n_0_2841), .B2(
      n_0_2778), .C1(n_0_2839), .C2(n_0_2747), .ZN(n_0_117_3));
   INV_X1 i_0_117_7 (.A(n_0_117_3), .ZN(n_0_2844));
   AOI222_X1 i_0_117_8 (.A1(n_0_2840), .A2(n_0_2811), .B1(n_0_2841), .B2(
      n_0_2779), .C1(n_0_2839), .C2(n_0_2748), .ZN(n_0_117_4));
   INV_X1 i_0_117_9 (.A(n_0_117_4), .ZN(n_0_2845));
   AOI222_X1 i_0_117_10 (.A1(n_0_2840), .A2(n_0_2812), .B1(n_0_2841), .B2(
      n_0_2780), .C1(n_0_2839), .C2(n_0_2749), .ZN(n_0_117_5));
   INV_X1 i_0_117_11 (.A(n_0_117_5), .ZN(n_0_2846));
   AOI222_X1 i_0_117_12 (.A1(n_0_2840), .A2(n_0_2813), .B1(n_0_2841), .B2(
      n_0_2781), .C1(n_0_2839), .C2(n_0_2750), .ZN(n_0_117_6));
   INV_X1 i_0_117_13 (.A(n_0_117_6), .ZN(n_0_2847));
   AOI222_X1 i_0_117_14 (.A1(n_0_2840), .A2(n_0_2814), .B1(n_0_2841), .B2(
      n_0_2782), .C1(n_0_2839), .C2(n_0_2751), .ZN(n_0_117_7));
   INV_X1 i_0_117_15 (.A(n_0_117_7), .ZN(n_0_2848));
   AOI222_X1 i_0_117_16 (.A1(n_0_2840), .A2(n_0_2815), .B1(n_0_2841), .B2(
      n_0_2783), .C1(n_0_2839), .C2(n_0_2752), .ZN(n_0_117_8));
   INV_X1 i_0_117_17 (.A(n_0_117_8), .ZN(n_0_2849));
   AOI222_X1 i_0_117_18 (.A1(n_0_2840), .A2(n_0_2816), .B1(n_0_2841), .B2(
      n_0_2784), .C1(n_0_2839), .C2(n_0_2753), .ZN(n_0_117_9));
   INV_X1 i_0_117_19 (.A(n_0_117_9), .ZN(n_0_2850));
   AOI222_X1 i_0_117_20 (.A1(n_0_2840), .A2(n_0_2817), .B1(n_0_2841), .B2(
      n_0_2785), .C1(n_0_2839), .C2(n_0_2754), .ZN(n_0_117_10));
   INV_X1 i_0_117_21 (.A(n_0_117_10), .ZN(n_0_2851));
   AOI222_X1 i_0_117_22 (.A1(n_0_2840), .A2(n_0_2818), .B1(n_0_2841), .B2(
      n_0_2786), .C1(n_0_2839), .C2(n_0_2755), .ZN(n_0_117_11));
   INV_X1 i_0_117_23 (.A(n_0_117_11), .ZN(n_0_2852));
   AOI222_X1 i_0_117_24 (.A1(n_0_2840), .A2(n_0_2819), .B1(n_0_2841), .B2(
      n_0_2787), .C1(n_0_2839), .C2(n_0_2756), .ZN(n_0_117_12));
   INV_X1 i_0_117_25 (.A(n_0_117_12), .ZN(n_0_2853));
   AOI222_X1 i_0_117_26 (.A1(n_0_2840), .A2(n_0_2820), .B1(n_0_2841), .B2(
      n_0_2788), .C1(n_0_2839), .C2(n_0_2757), .ZN(n_0_117_13));
   INV_X1 i_0_117_27 (.A(n_0_117_13), .ZN(n_0_2854));
   AOI222_X1 i_0_117_28 (.A1(n_0_2840), .A2(n_0_2821), .B1(n_0_2841), .B2(
      n_0_2789), .C1(n_0_2839), .C2(n_0_2758), .ZN(n_0_117_14));
   INV_X1 i_0_117_29 (.A(n_0_117_14), .ZN(n_0_2855));
   AOI222_X1 i_0_117_30 (.A1(n_0_2840), .A2(n_0_2822), .B1(n_0_2841), .B2(
      n_0_2790), .C1(n_0_2839), .C2(n_0_2759), .ZN(n_0_117_15));
   INV_X1 i_0_117_31 (.A(n_0_117_15), .ZN(n_0_2856));
   AOI222_X1 i_0_117_32 (.A1(n_0_2840), .A2(n_0_2823), .B1(n_0_2841), .B2(
      n_0_2791), .C1(n_0_2839), .C2(n_0_2760), .ZN(n_0_117_16));
   INV_X1 i_0_117_33 (.A(n_0_117_16), .ZN(n_0_2857));
   AOI222_X1 i_0_117_34 (.A1(n_0_2840), .A2(n_0_2824), .B1(n_0_2841), .B2(
      n_0_2792), .C1(n_0_2839), .C2(n_0_2761), .ZN(n_0_117_17));
   INV_X1 i_0_117_35 (.A(n_0_117_17), .ZN(n_0_2858));
   AOI222_X1 i_0_117_36 (.A1(n_0_2840), .A2(n_0_2825), .B1(n_0_2841), .B2(
      n_0_2793), .C1(n_0_2839), .C2(n_0_2762), .ZN(n_0_117_18));
   INV_X1 i_0_117_37 (.A(n_0_117_18), .ZN(n_0_2859));
   AOI222_X1 i_0_117_38 (.A1(n_0_2840), .A2(n_0_2826), .B1(n_0_2841), .B2(
      n_0_2794), .C1(n_0_2839), .C2(n_0_2763), .ZN(n_0_117_19));
   INV_X1 i_0_117_39 (.A(n_0_117_19), .ZN(n_0_2860));
   AOI222_X1 i_0_117_40 (.A1(n_0_2840), .A2(n_0_2827), .B1(n_0_2841), .B2(
      n_0_2795), .C1(n_0_2839), .C2(n_0_2764), .ZN(n_0_117_20));
   INV_X1 i_0_117_41 (.A(n_0_117_20), .ZN(n_0_2861));
   AOI222_X1 i_0_117_42 (.A1(n_0_2840), .A2(n_0_2828), .B1(n_0_2841), .B2(
      n_0_2796), .C1(n_0_2839), .C2(n_0_2765), .ZN(n_0_117_21));
   INV_X1 i_0_117_43 (.A(n_0_117_21), .ZN(n_0_2862));
   AOI222_X1 i_0_117_44 (.A1(n_0_2840), .A2(n_0_2829), .B1(n_0_2841), .B2(
      n_0_2797), .C1(n_0_2839), .C2(n_0_2766), .ZN(n_0_117_22));
   INV_X1 i_0_117_45 (.A(n_0_117_22), .ZN(n_0_2863));
   AOI222_X1 i_0_117_46 (.A1(n_0_2840), .A2(n_0_2830), .B1(n_0_2841), .B2(
      n_0_2798), .C1(n_0_2839), .C2(n_0_2767), .ZN(n_0_117_23));
   INV_X1 i_0_117_47 (.A(n_0_117_23), .ZN(n_0_2864));
   AOI222_X1 i_0_117_48 (.A1(n_0_2840), .A2(n_0_2831), .B1(n_0_2841), .B2(
      n_0_2799), .C1(n_0_2839), .C2(n_0_2768), .ZN(n_0_117_24));
   INV_X1 i_0_117_49 (.A(n_0_117_24), .ZN(n_0_2865));
   AOI222_X1 i_0_117_50 (.A1(n_0_2840), .A2(n_0_2832), .B1(n_0_2841), .B2(
      n_0_2800), .C1(n_0_2839), .C2(n_0_2769), .ZN(n_0_117_25));
   INV_X1 i_0_117_51 (.A(n_0_117_25), .ZN(n_0_2866));
   AOI222_X1 i_0_117_52 (.A1(n_0_2840), .A2(n_0_2833), .B1(n_0_2841), .B2(
      n_0_2801), .C1(n_0_2839), .C2(n_0_2770), .ZN(n_0_117_26));
   INV_X1 i_0_117_53 (.A(n_0_117_26), .ZN(n_0_2867));
   AOI222_X1 i_0_117_54 (.A1(n_0_2840), .A2(n_0_2834), .B1(n_0_2841), .B2(
      n_0_2802), .C1(n_0_2839), .C2(n_0_2771), .ZN(n_0_117_27));
   INV_X1 i_0_117_55 (.A(n_0_117_27), .ZN(n_0_2868));
   AOI222_X1 i_0_117_56 (.A1(n_0_2840), .A2(n_0_2835), .B1(n_0_2841), .B2(
      n_0_2803), .C1(n_0_2839), .C2(n_0_2772), .ZN(n_0_117_28));
   INV_X1 i_0_117_57 (.A(n_0_117_28), .ZN(n_0_2869));
   AOI222_X1 i_0_117_58 (.A1(n_0_2840), .A2(n_0_2836), .B1(n_0_2841), .B2(
      n_0_2804), .C1(n_0_2839), .C2(n_0_2773), .ZN(n_0_117_29));
   INV_X1 i_0_117_59 (.A(n_0_117_29), .ZN(n_0_2870));
   AND2_X1 i_0_117_60 (.A1(n_0_2839), .A2(n_0_2774), .ZN(n_0_117_30));
   AOI221_X1 i_0_117_61 (.A(n_0_117_30), .B1(n_0_2840), .B2(n_0_2837), .C1(
      n_0_2841), .C2(n_0_2805), .ZN(n_0_117_31));
   INV_X1 i_0_117_62 (.A(n_0_117_31), .ZN(n_0_2871));
   AOI221_X1 i_0_117_63 (.A(n_0_117_30), .B1(n_0_2840), .B2(n_0_2838), .C1(
      n_0_2841), .C2(n_0_2806), .ZN(n_0_117_32));
   INV_X1 i_0_117_64 (.A(n_0_117_32), .ZN(n_0_2872));
   datapath__0_116 i_0_118 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_59, 
      n_0_2872, n_0_2871, n_0_2870, n_0_2869, n_0_2868, n_0_2867, n_0_2866, 
      n_0_2865, n_0_2864, n_0_2863, n_0_2862, n_0_2861, n_0_2860, n_0_2859, 
      n_0_2858, n_0_2857, n_0_2856, n_0_2855, n_0_2854, n_0_2853, n_0_2852, 
      n_0_2851, n_0_2850, n_0_2849, n_0_2848, n_0_2847, n_0_2846, n_0_2845, 
      n_0_2844, n_0_2843, n_0_2842}), .p_2({n_0_2904, n_0_2903, n_0_2902, 
      n_0_2901, n_0_2900, n_0_2899, n_0_2898, n_0_2897, n_0_2896, n_0_2895, 
      n_0_2894, n_0_2893, n_0_2892, n_0_2891, n_0_2890, n_0_2889, n_0_2888, 
      n_0_2887, n_0_2886, n_0_2885, n_0_2884, n_0_2883, n_0_2882, n_0_2881, 
      n_0_2880, n_0_2879, n_0_2878, n_0_2877, n_0_2876, n_0_2875, n_0_2874, 
      n_0_2873}));
   datapath__0_117 i_0_119 (.multiplicand2(multiplicand2), .p_0({uc_60, n_0_2872, 
      n_0_2871, n_0_2870, n_0_2869, n_0_2868, n_0_2867, n_0_2866, n_0_2865, 
      n_0_2864, n_0_2863, n_0_2862, n_0_2861, n_0_2860, n_0_2859, n_0_2858, 
      n_0_2857, n_0_2856, n_0_2855, n_0_2854, n_0_2853, n_0_2852, n_0_2851, 
      n_0_2850, n_0_2849, n_0_2848, n_0_2847, n_0_2846, n_0_2845, n_0_2844, 
      n_0_2843, n_0_2842}), .p_1({n_0_2936, n_0_2935, n_0_2934, n_0_2933, 
      n_0_2932, n_0_2931, n_0_2930, n_0_2929, n_0_2928, n_0_2927, n_0_2926, 
      n_0_2925, n_0_2924, n_0_2923, n_0_2922, n_0_2921, n_0_2920, n_0_2919, 
      n_0_2918, n_0_2917, n_0_2916, n_0_2915, n_0_2914, n_0_2913, n_0_2912, 
      n_0_2911, n_0_2910, n_0_2909, n_0_2908, n_0_2907, n_0_2906, n_0_2905}));
   INV_X1 i_0_120_0 (.A(multiplier2[30]), .ZN(n_0_120_0));
   AND2_X1 i_0_120_1 (.A1(n_0_120_0), .A2(multiplier2[29]), .ZN(n_0_2938));
   NOR2_X1 i_0_120_2 (.A1(n_0_120_0), .A2(multiplier2[29]), .ZN(n_0_2939));
   NOR2_X1 i_0_120_3 (.A1(n_0_2938), .A2(n_0_2939), .ZN(n_0_2937));
   AOI222_X1 i_0_121_0 (.A1(n_0_2905), .A2(n_0_2938), .B1(n_0_2873), .B2(
      n_0_2939), .C1(n_0_2842), .C2(n_0_2937), .ZN(n_0_121_0));
   INV_X1 i_0_121_1 (.A(n_0_121_0), .ZN(product[30]));
   AOI222_X1 i_0_121_2 (.A1(n_0_2938), .A2(n_0_2906), .B1(n_0_2939), .B2(
      n_0_2874), .C1(n_0_2937), .C2(n_0_2843), .ZN(n_0_121_1));
   INV_X1 i_0_121_3 (.A(n_0_121_1), .ZN(n_0_2940));
   AOI222_X1 i_0_121_4 (.A1(n_0_2938), .A2(n_0_2907), .B1(n_0_2939), .B2(
      n_0_2875), .C1(n_0_2937), .C2(n_0_2844), .ZN(n_0_121_2));
   INV_X1 i_0_121_5 (.A(n_0_121_2), .ZN(n_0_2941));
   AOI222_X1 i_0_121_6 (.A1(n_0_2938), .A2(n_0_2908), .B1(n_0_2939), .B2(
      n_0_2876), .C1(n_0_2937), .C2(n_0_2845), .ZN(n_0_121_3));
   INV_X1 i_0_121_7 (.A(n_0_121_3), .ZN(n_0_2942));
   AOI222_X1 i_0_121_8 (.A1(n_0_2938), .A2(n_0_2909), .B1(n_0_2939), .B2(
      n_0_2877), .C1(n_0_2937), .C2(n_0_2846), .ZN(n_0_121_4));
   INV_X1 i_0_121_9 (.A(n_0_121_4), .ZN(n_0_2943));
   AOI222_X1 i_0_121_10 (.A1(n_0_2938), .A2(n_0_2910), .B1(n_0_2939), .B2(
      n_0_2878), .C1(n_0_2937), .C2(n_0_2847), .ZN(n_0_121_5));
   INV_X1 i_0_121_11 (.A(n_0_121_5), .ZN(n_0_2944));
   AOI222_X1 i_0_121_12 (.A1(n_0_2938), .A2(n_0_2911), .B1(n_0_2939), .B2(
      n_0_2879), .C1(n_0_2937), .C2(n_0_2848), .ZN(n_0_121_6));
   INV_X1 i_0_121_13 (.A(n_0_121_6), .ZN(n_0_2945));
   AOI222_X1 i_0_121_14 (.A1(n_0_2938), .A2(n_0_2912), .B1(n_0_2939), .B2(
      n_0_2880), .C1(n_0_2937), .C2(n_0_2849), .ZN(n_0_121_7));
   INV_X1 i_0_121_15 (.A(n_0_121_7), .ZN(n_0_2946));
   AOI222_X1 i_0_121_16 (.A1(n_0_2938), .A2(n_0_2913), .B1(n_0_2939), .B2(
      n_0_2881), .C1(n_0_2937), .C2(n_0_2850), .ZN(n_0_121_8));
   INV_X1 i_0_121_17 (.A(n_0_121_8), .ZN(n_0_2947));
   AOI222_X1 i_0_121_18 (.A1(n_0_2938), .A2(n_0_2914), .B1(n_0_2939), .B2(
      n_0_2882), .C1(n_0_2937), .C2(n_0_2851), .ZN(n_0_121_9));
   INV_X1 i_0_121_19 (.A(n_0_121_9), .ZN(n_0_2948));
   AOI222_X1 i_0_121_20 (.A1(n_0_2938), .A2(n_0_2915), .B1(n_0_2939), .B2(
      n_0_2883), .C1(n_0_2937), .C2(n_0_2852), .ZN(n_0_121_10));
   INV_X1 i_0_121_21 (.A(n_0_121_10), .ZN(n_0_2949));
   AOI222_X1 i_0_121_22 (.A1(n_0_2938), .A2(n_0_2916), .B1(n_0_2939), .B2(
      n_0_2884), .C1(n_0_2937), .C2(n_0_2853), .ZN(n_0_121_11));
   INV_X1 i_0_121_23 (.A(n_0_121_11), .ZN(n_0_2950));
   AOI222_X1 i_0_121_24 (.A1(n_0_2938), .A2(n_0_2917), .B1(n_0_2939), .B2(
      n_0_2885), .C1(n_0_2937), .C2(n_0_2854), .ZN(n_0_121_12));
   INV_X1 i_0_121_25 (.A(n_0_121_12), .ZN(n_0_2951));
   AOI222_X1 i_0_121_26 (.A1(n_0_2938), .A2(n_0_2918), .B1(n_0_2939), .B2(
      n_0_2886), .C1(n_0_2937), .C2(n_0_2855), .ZN(n_0_121_13));
   INV_X1 i_0_121_27 (.A(n_0_121_13), .ZN(n_0_2952));
   AOI222_X1 i_0_121_28 (.A1(n_0_2938), .A2(n_0_2919), .B1(n_0_2939), .B2(
      n_0_2887), .C1(n_0_2937), .C2(n_0_2856), .ZN(n_0_121_14));
   INV_X1 i_0_121_29 (.A(n_0_121_14), .ZN(n_0_2953));
   AOI222_X1 i_0_121_30 (.A1(n_0_2938), .A2(n_0_2920), .B1(n_0_2939), .B2(
      n_0_2888), .C1(n_0_2937), .C2(n_0_2857), .ZN(n_0_121_15));
   INV_X1 i_0_121_31 (.A(n_0_121_15), .ZN(n_0_2954));
   AOI222_X1 i_0_121_32 (.A1(n_0_2938), .A2(n_0_2921), .B1(n_0_2939), .B2(
      n_0_2889), .C1(n_0_2937), .C2(n_0_2858), .ZN(n_0_121_16));
   INV_X1 i_0_121_33 (.A(n_0_121_16), .ZN(n_0_2955));
   AOI222_X1 i_0_121_34 (.A1(n_0_2938), .A2(n_0_2922), .B1(n_0_2939), .B2(
      n_0_2890), .C1(n_0_2937), .C2(n_0_2859), .ZN(n_0_121_17));
   INV_X1 i_0_121_35 (.A(n_0_121_17), .ZN(n_0_2956));
   AOI222_X1 i_0_121_36 (.A1(n_0_2938), .A2(n_0_2923), .B1(n_0_2939), .B2(
      n_0_2891), .C1(n_0_2937), .C2(n_0_2860), .ZN(n_0_121_18));
   INV_X1 i_0_121_37 (.A(n_0_121_18), .ZN(n_0_2957));
   AOI222_X1 i_0_121_38 (.A1(n_0_2938), .A2(n_0_2924), .B1(n_0_2939), .B2(
      n_0_2892), .C1(n_0_2937), .C2(n_0_2861), .ZN(n_0_121_19));
   INV_X1 i_0_121_39 (.A(n_0_121_19), .ZN(n_0_2958));
   AOI222_X1 i_0_121_40 (.A1(n_0_2938), .A2(n_0_2925), .B1(n_0_2939), .B2(
      n_0_2893), .C1(n_0_2937), .C2(n_0_2862), .ZN(n_0_121_20));
   INV_X1 i_0_121_41 (.A(n_0_121_20), .ZN(n_0_2959));
   AOI222_X1 i_0_121_42 (.A1(n_0_2938), .A2(n_0_2926), .B1(n_0_2939), .B2(
      n_0_2894), .C1(n_0_2937), .C2(n_0_2863), .ZN(n_0_121_21));
   INV_X1 i_0_121_43 (.A(n_0_121_21), .ZN(n_0_2960));
   AOI222_X1 i_0_121_44 (.A1(n_0_2938), .A2(n_0_2927), .B1(n_0_2939), .B2(
      n_0_2895), .C1(n_0_2937), .C2(n_0_2864), .ZN(n_0_121_22));
   INV_X1 i_0_121_45 (.A(n_0_121_22), .ZN(n_0_2961));
   AOI222_X1 i_0_121_46 (.A1(n_0_2938), .A2(n_0_2928), .B1(n_0_2939), .B2(
      n_0_2896), .C1(n_0_2937), .C2(n_0_2865), .ZN(n_0_121_23));
   INV_X1 i_0_121_47 (.A(n_0_121_23), .ZN(n_0_2962));
   AOI222_X1 i_0_121_48 (.A1(n_0_2938), .A2(n_0_2929), .B1(n_0_2939), .B2(
      n_0_2897), .C1(n_0_2937), .C2(n_0_2866), .ZN(n_0_121_24));
   INV_X1 i_0_121_49 (.A(n_0_121_24), .ZN(n_0_2963));
   AOI222_X1 i_0_121_50 (.A1(n_0_2938), .A2(n_0_2930), .B1(n_0_2939), .B2(
      n_0_2898), .C1(n_0_2937), .C2(n_0_2867), .ZN(n_0_121_25));
   INV_X1 i_0_121_51 (.A(n_0_121_25), .ZN(n_0_2964));
   AOI222_X1 i_0_121_52 (.A1(n_0_2938), .A2(n_0_2931), .B1(n_0_2939), .B2(
      n_0_2899), .C1(n_0_2937), .C2(n_0_2868), .ZN(n_0_121_26));
   INV_X1 i_0_121_53 (.A(n_0_121_26), .ZN(n_0_2965));
   AOI222_X1 i_0_121_54 (.A1(n_0_2938), .A2(n_0_2932), .B1(n_0_2939), .B2(
      n_0_2900), .C1(n_0_2937), .C2(n_0_2869), .ZN(n_0_121_27));
   INV_X1 i_0_121_55 (.A(n_0_121_27), .ZN(n_0_2966));
   AOI222_X1 i_0_121_56 (.A1(n_0_2938), .A2(n_0_2933), .B1(n_0_2939), .B2(
      n_0_2901), .C1(n_0_2937), .C2(n_0_2870), .ZN(n_0_121_28));
   INV_X1 i_0_121_57 (.A(n_0_121_28), .ZN(n_0_2967));
   AOI222_X1 i_0_121_58 (.A1(n_0_2938), .A2(n_0_2934), .B1(n_0_2939), .B2(
      n_0_2902), .C1(n_0_2937), .C2(n_0_2871), .ZN(n_0_121_29));
   INV_X1 i_0_121_59 (.A(n_0_121_29), .ZN(n_0_2968));
   AND2_X1 i_0_121_60 (.A1(n_0_2937), .A2(n_0_2872), .ZN(n_0_121_30));
   AOI221_X1 i_0_121_61 (.A(n_0_121_30), .B1(n_0_2938), .B2(n_0_2935), .C1(
      n_0_2939), .C2(n_0_2903), .ZN(n_0_121_31));
   INV_X1 i_0_121_62 (.A(n_0_121_31), .ZN(n_0_2969));
   AOI221_X1 i_0_121_63 (.A(n_0_121_30), .B1(n_0_2938), .B2(n_0_2936), .C1(
      n_0_2939), .C2(n_0_2904), .ZN(n_0_121_32));
   INV_X1 i_0_121_64 (.A(n_0_121_32), .ZN(n_0_2970));
   datapath__0_120 i_0_122 (.p_0({n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, multiplicand2[0]}), .p_1({uc_61, 
      n_0_2970, n_0_2969, n_0_2968, n_0_2967, n_0_2966, n_0_2965, n_0_2964, 
      n_0_2963, n_0_2962, n_0_2961, n_0_2960, n_0_2959, n_0_2958, n_0_2957, 
      n_0_2956, n_0_2955, n_0_2954, n_0_2953, n_0_2952, n_0_2951, n_0_2950, 
      n_0_2949, n_0_2948, n_0_2947, n_0_2946, n_0_2945, n_0_2944, n_0_2943, 
      n_0_2942, n_0_2941, n_0_2940}), .p_2({n_0_3002, n_0_3001, n_0_3000, 
      n_0_2999, n_0_2998, n_0_2997, n_0_2996, n_0_2995, n_0_2994, n_0_2993, 
      n_0_2992, n_0_2991, n_0_2990, n_0_2989, n_0_2988, n_0_2987, n_0_2986, 
      n_0_2985, n_0_2984, n_0_2983, n_0_2982, n_0_2981, n_0_2980, n_0_2979, 
      n_0_2978, n_0_2977, n_0_2976, n_0_2975, n_0_2974, n_0_2973, n_0_2972, 
      n_0_2971}));
   datapath__0_121 i_0_123 (.multiplicand2(multiplicand2), .p_0({uc_62, n_0_2970, 
      n_0_2969, n_0_2968, n_0_2967, n_0_2966, n_0_2965, n_0_2964, n_0_2963, 
      n_0_2962, n_0_2961, n_0_2960, n_0_2959, n_0_2958, n_0_2957, n_0_2956, 
      n_0_2955, n_0_2954, n_0_2953, n_0_2952, n_0_2951, n_0_2950, n_0_2949, 
      n_0_2948, n_0_2947, n_0_2946, n_0_2945, n_0_2944, n_0_2943, n_0_2942, 
      n_0_2941, n_0_2940}), .p_1({n_0_3034, n_0_3033, n_0_3032, n_0_3031, 
      n_0_3030, n_0_3029, n_0_3028, n_0_3027, n_0_3026, n_0_3025, n_0_3024, 
      n_0_3023, n_0_3022, n_0_3021, n_0_3020, n_0_3019, n_0_3018, n_0_3017, 
      n_0_3016, n_0_3015, n_0_3014, n_0_3013, n_0_3012, n_0_3011, n_0_3010, 
      n_0_3009, n_0_3008, n_0_3007, n_0_3006, n_0_3005, n_0_3004, n_0_3003}));
   INV_X1 i_0_124_0 (.A(multiplier2[31]), .ZN(n_0_124_0));
   AND2_X1 i_0_124_1 (.A1(n_0_124_0), .A2(multiplier2[30]), .ZN(n_0_3036));
   NOR2_X1 i_0_124_2 (.A1(n_0_124_0), .A2(multiplier2[30]), .ZN(n_0_3037));
   NOR2_X1 i_0_124_3 (.A1(n_0_3036), .A2(n_0_3037), .ZN(n_0_3035));
   AOI222_X1 i_0_125_0 (.A1(n_0_3003), .A2(n_0_3036), .B1(n_0_2971), .B2(
      n_0_3037), .C1(n_0_2940), .C2(n_0_3035), .ZN(n_0_125_0));
   INV_X1 i_0_125_1 (.A(n_0_125_0), .ZN(product[31]));
   AOI222_X1 i_0_125_2 (.A1(n_0_3036), .A2(n_0_3004), .B1(n_0_3037), .B2(
      n_0_2972), .C1(n_0_3035), .C2(n_0_2941), .ZN(n_0_125_1));
   INV_X1 i_0_125_3 (.A(n_0_125_1), .ZN(product[32]));
   AOI222_X1 i_0_125_4 (.A1(n_0_3036), .A2(n_0_3005), .B1(n_0_3037), .B2(
      n_0_2973), .C1(n_0_3035), .C2(n_0_2942), .ZN(n_0_125_2));
   INV_X1 i_0_125_5 (.A(n_0_125_2), .ZN(product[33]));
   AOI222_X1 i_0_125_6 (.A1(n_0_3036), .A2(n_0_3006), .B1(n_0_3037), .B2(
      n_0_2974), .C1(n_0_3035), .C2(n_0_2943), .ZN(n_0_125_3));
   INV_X1 i_0_125_7 (.A(n_0_125_3), .ZN(product[34]));
   AOI222_X1 i_0_125_8 (.A1(n_0_3036), .A2(n_0_3007), .B1(n_0_3037), .B2(
      n_0_2975), .C1(n_0_3035), .C2(n_0_2944), .ZN(n_0_125_4));
   INV_X1 i_0_125_9 (.A(n_0_125_4), .ZN(product[35]));
   AOI222_X1 i_0_125_10 (.A1(n_0_3036), .A2(n_0_3008), .B1(n_0_3037), .B2(
      n_0_2976), .C1(n_0_3035), .C2(n_0_2945), .ZN(n_0_125_5));
   INV_X1 i_0_125_11 (.A(n_0_125_5), .ZN(product[36]));
   AOI222_X1 i_0_125_12 (.A1(n_0_3036), .A2(n_0_3009), .B1(n_0_3037), .B2(
      n_0_2977), .C1(n_0_3035), .C2(n_0_2946), .ZN(n_0_125_6));
   INV_X1 i_0_125_13 (.A(n_0_125_6), .ZN(product[37]));
   AOI222_X1 i_0_125_14 (.A1(n_0_3036), .A2(n_0_3010), .B1(n_0_3037), .B2(
      n_0_2978), .C1(n_0_3035), .C2(n_0_2947), .ZN(n_0_125_7));
   INV_X1 i_0_125_15 (.A(n_0_125_7), .ZN(product[38]));
   AOI222_X1 i_0_125_16 (.A1(n_0_3036), .A2(n_0_3011), .B1(n_0_3037), .B2(
      n_0_2979), .C1(n_0_3035), .C2(n_0_2948), .ZN(n_0_125_8));
   INV_X1 i_0_125_17 (.A(n_0_125_8), .ZN(product[39]));
   AOI222_X1 i_0_125_18 (.A1(n_0_3036), .A2(n_0_3012), .B1(n_0_3037), .B2(
      n_0_2980), .C1(n_0_3035), .C2(n_0_2949), .ZN(n_0_125_9));
   INV_X1 i_0_125_19 (.A(n_0_125_9), .ZN(product[40]));
   AOI222_X1 i_0_125_20 (.A1(n_0_3036), .A2(n_0_3013), .B1(n_0_3037), .B2(
      n_0_2981), .C1(n_0_3035), .C2(n_0_2950), .ZN(n_0_125_10));
   INV_X1 i_0_125_21 (.A(n_0_125_10), .ZN(product[41]));
   AOI222_X1 i_0_125_22 (.A1(n_0_3036), .A2(n_0_3014), .B1(n_0_3037), .B2(
      n_0_2982), .C1(n_0_3035), .C2(n_0_2951), .ZN(n_0_125_11));
   INV_X1 i_0_125_23 (.A(n_0_125_11), .ZN(product[42]));
   AOI222_X1 i_0_125_24 (.A1(n_0_3036), .A2(n_0_3015), .B1(n_0_3037), .B2(
      n_0_2983), .C1(n_0_3035), .C2(n_0_2952), .ZN(n_0_125_12));
   INV_X1 i_0_125_25 (.A(n_0_125_12), .ZN(product[43]));
   AOI222_X1 i_0_125_26 (.A1(n_0_3036), .A2(n_0_3016), .B1(n_0_3037), .B2(
      n_0_2984), .C1(n_0_3035), .C2(n_0_2953), .ZN(n_0_125_13));
   INV_X1 i_0_125_27 (.A(n_0_125_13), .ZN(product[44]));
   AOI222_X1 i_0_125_28 (.A1(n_0_3036), .A2(n_0_3017), .B1(n_0_3037), .B2(
      n_0_2985), .C1(n_0_3035), .C2(n_0_2954), .ZN(n_0_125_14));
   INV_X1 i_0_125_29 (.A(n_0_125_14), .ZN(product[45]));
   AOI222_X1 i_0_125_30 (.A1(n_0_3036), .A2(n_0_3018), .B1(n_0_3037), .B2(
      n_0_2986), .C1(n_0_3035), .C2(n_0_2955), .ZN(n_0_125_15));
   INV_X1 i_0_125_31 (.A(n_0_125_15), .ZN(product[46]));
   AOI222_X1 i_0_125_32 (.A1(n_0_3036), .A2(n_0_3019), .B1(n_0_3037), .B2(
      n_0_2987), .C1(n_0_3035), .C2(n_0_2956), .ZN(n_0_125_16));
   INV_X1 i_0_125_33 (.A(n_0_125_16), .ZN(product[47]));
   AOI222_X1 i_0_125_34 (.A1(n_0_3036), .A2(n_0_3020), .B1(n_0_3037), .B2(
      n_0_2988), .C1(n_0_3035), .C2(n_0_2957), .ZN(n_0_125_17));
   INV_X1 i_0_125_35 (.A(n_0_125_17), .ZN(product[48]));
   AOI222_X1 i_0_125_36 (.A1(n_0_3036), .A2(n_0_3021), .B1(n_0_3037), .B2(
      n_0_2989), .C1(n_0_3035), .C2(n_0_2958), .ZN(n_0_125_18));
   INV_X1 i_0_125_37 (.A(n_0_125_18), .ZN(product[49]));
   AOI222_X1 i_0_125_38 (.A1(n_0_3036), .A2(n_0_3022), .B1(n_0_3037), .B2(
      n_0_2990), .C1(n_0_3035), .C2(n_0_2959), .ZN(n_0_125_19));
   INV_X1 i_0_125_39 (.A(n_0_125_19), .ZN(product[50]));
   AOI222_X1 i_0_125_40 (.A1(n_0_3036), .A2(n_0_3023), .B1(n_0_3037), .B2(
      n_0_2991), .C1(n_0_3035), .C2(n_0_2960), .ZN(n_0_125_20));
   INV_X1 i_0_125_41 (.A(n_0_125_20), .ZN(product[51]));
   AOI222_X1 i_0_125_42 (.A1(n_0_3036), .A2(n_0_3024), .B1(n_0_3037), .B2(
      n_0_2992), .C1(n_0_3035), .C2(n_0_2961), .ZN(n_0_125_21));
   INV_X1 i_0_125_43 (.A(n_0_125_21), .ZN(product[52]));
   AOI222_X1 i_0_125_44 (.A1(n_0_3036), .A2(n_0_3025), .B1(n_0_3037), .B2(
      n_0_2993), .C1(n_0_3035), .C2(n_0_2962), .ZN(n_0_125_22));
   INV_X1 i_0_125_45 (.A(n_0_125_22), .ZN(product[53]));
   AOI222_X1 i_0_125_46 (.A1(n_0_3036), .A2(n_0_3026), .B1(n_0_3037), .B2(
      n_0_2994), .C1(n_0_3035), .C2(n_0_2963), .ZN(n_0_125_23));
   INV_X1 i_0_125_47 (.A(n_0_125_23), .ZN(product[54]));
   AOI222_X1 i_0_125_48 (.A1(n_0_3036), .A2(n_0_3027), .B1(n_0_3037), .B2(
      n_0_2995), .C1(n_0_3035), .C2(n_0_2964), .ZN(n_0_125_24));
   INV_X1 i_0_125_49 (.A(n_0_125_24), .ZN(product[55]));
   AOI222_X1 i_0_125_50 (.A1(n_0_3036), .A2(n_0_3028), .B1(n_0_3037), .B2(
      n_0_2996), .C1(n_0_3035), .C2(n_0_2965), .ZN(n_0_125_25));
   INV_X1 i_0_125_51 (.A(n_0_125_25), .ZN(product[56]));
   AOI222_X1 i_0_125_52 (.A1(n_0_3036), .A2(n_0_3029), .B1(n_0_3037), .B2(
      n_0_2997), .C1(n_0_3035), .C2(n_0_2966), .ZN(n_0_125_26));
   INV_X1 i_0_125_53 (.A(n_0_125_26), .ZN(product[57]));
   AOI222_X1 i_0_125_54 (.A1(n_0_3036), .A2(n_0_3030), .B1(n_0_3037), .B2(
      n_0_2998), .C1(n_0_3035), .C2(n_0_2967), .ZN(n_0_125_27));
   INV_X1 i_0_125_55 (.A(n_0_125_27), .ZN(product[58]));
   AOI222_X1 i_0_125_56 (.A1(n_0_3036), .A2(n_0_3031), .B1(n_0_3037), .B2(
      n_0_2999), .C1(n_0_3035), .C2(n_0_2968), .ZN(n_0_125_28));
   INV_X1 i_0_125_57 (.A(n_0_125_28), .ZN(product[59]));
   AOI222_X1 i_0_125_58 (.A1(n_0_3036), .A2(n_0_3032), .B1(n_0_3037), .B2(
      n_0_3000), .C1(n_0_3035), .C2(n_0_2969), .ZN(n_0_125_29));
   INV_X1 i_0_125_59 (.A(n_0_125_29), .ZN(product[60]));
   AND2_X1 i_0_125_60 (.A1(n_0_3035), .A2(n_0_2970), .ZN(n_0_125_30));
   AOI221_X1 i_0_125_61 (.A(n_0_125_30), .B1(n_0_3036), .B2(n_0_3033), .C1(
      n_0_3037), .C2(n_0_3001), .ZN(n_0_125_31));
   INV_X1 i_0_125_62 (.A(n_0_125_31), .ZN(product[61]));
   AOI221_X1 i_0_125_63 (.A(n_0_125_30), .B1(n_0_3036), .B2(n_0_3034), .C1(
      n_0_3037), .C2(n_0_3002), .ZN(n_0_125_32));
   INV_X1 i_0_125_64 (.A(n_0_125_32), .ZN(product[62]));
endmodule

module boothMult(i_clk, i_rst, i_en, i_inputA, i_inputB, o_result);
   input i_clk;
   input i_rst;
   input i_en;
   input [31:0]i_inputA;
   input [31:0]i_inputB;
   output [63:0]o_result;

   wire [31:0]B_reg;
   wire [31:0]A_reg;
   wire [63:0]out_reg;

   registerNbits_bbox_0 regB (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(
      i_inputB), .p_4(B_reg));
   registerNbits_bbox_1 outReg (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(
      out_reg), .p_4(o_result));
   registerNbits_bbox regA (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(i_inputA), 
      .p_4(A_reg));
   booth boothUnit (.multiplicand2(A_reg), .multiplier2(B_reg), .product(out_reg));
endmodule
