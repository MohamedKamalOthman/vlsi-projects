module HA (
	input a,
	input b,
	output sum,
	output carry
);
assign {carry, sum} = a + b;
endmodule

module FA (
	input a,
	input b,
	input c,
	output sum,
	output carry
);
assign {carry, sum} = a + b + c;
endmodule

module signed_wallace_tree_multipler #(parameter SIZE = 32)(
	input [SIZE - 1:0] A,
	input [SIZE - 1:0] B,
	output [2 * SIZE - 1:0] result
);
reg [SIZE - 1:0] p[SIZE - 1:0];
// Set First 32 x 32 Products Of A x B
integer i;
always @(*) begin
	for(i = 0;i <= SIZE - 1;i = i + 1)begin
		if(i == SIZE - 1)  
			p[i] = {(A[i] & B[(SIZE - 1)]), ~({(SIZE - 1){A[i]}} & B[(SIZE - 2):0])};
		else
			p[i] = {~(A[i] & B[(SIZE - 1)]), {(SIZE - 1){A[i]}} & B[(SIZE - 2):0]};
	end
end

wire [1348:0] r;
wire [1348:0] c;

HA HA_0(p[0][1], p[1][0], r[0], c[0]);
FA FA_0(p[0][2], p[1][1], p[2][0], r[1], c[1]);
FA FA_1(p[0][3], p[1][2], p[2][1], r[2], c[2]);
HA HA_1(p[3][0], c[1], r[3], c[3]);
FA FA_2(p[0][4], p[1][3], p[2][2], r[4], c[4]);
FA FA_3(p[0][5], p[1][4], p[2][3], r[5], c[5]);
FA FA_4(p[0][6], p[1][5], p[2][4], r[6], c[6]);
HA HA_2(p[3][3], p[4][2], r[7], c[7]);
FA FA_5(p[0][7], p[1][6], p[2][5], r[8], c[8]);
FA FA_6(p[0][8], p[1][7], p[2][6], r[9], c[9]);
FA FA_7(p[0][9], p[1][8], p[2][7], r[10], c[10]);
HA HA_3(p[3][6], p[4][5], r[11], c[11]);
FA FA_8(p[0][10], p[1][9], p[2][8], r[12], c[12]);
FA FA_9(p[3][7], p[4][6], p[5][5], r[13], c[13]);
FA FA_10(p[0][11], p[1][10], p[2][9], r[14], c[14]);
FA FA_11(p[3][8], p[4][7], p[5][6], r[15], c[15]);
HA HA_4(p[6][5], p[7][4], r[16], c[16]);
FA FA_12(p[0][12], p[1][11], p[2][10], r[17], c[17]);
FA FA_13(p[3][9], p[4][8], p[5][7], r[18], c[18]);
FA FA_14(p[0][13], p[1][12], p[2][11], r[19], c[19]);
FA FA_15(p[3][10], p[4][9], p[5][8], r[20], c[20]);
FA FA_16(p[0][14], p[1][13], p[2][12], r[21], c[21]);
FA FA_17(p[3][11], p[4][10], p[5][9], r[22], c[22]);
HA HA_5(p[6][8], p[7][7], r[23], c[23]);
FA FA_18(p[0][15], p[1][14], p[2][13], r[24], c[24]);
FA FA_19(p[3][12], p[4][11], p[5][10], r[25], c[25]);
FA FA_20(p[0][16], p[1][15], p[2][14], r[26], c[26]);
FA FA_21(p[3][13], p[4][12], p[5][11], r[27], c[27]);
FA FA_22(p[0][17], p[1][16], p[2][15], r[28], c[28]);
FA FA_23(p[3][14], p[4][13], p[5][12], r[29], c[29]);
HA HA_6(p[6][11], p[7][10], r[30], c[30]);
FA FA_24(p[0][18], p[1][17], p[2][16], r[31], c[31]);
FA FA_25(p[3][15], p[4][14], p[5][13], r[32], c[32]);
FA FA_26(p[6][12], p[7][11], p[8][10], r[33], c[33]);
FA FA_27(p[0][19], p[1][18], p[2][17], r[34], c[34]);
FA FA_28(p[3][16], p[4][15], p[5][14], r[35], c[35]);
FA FA_29(p[6][13], p[7][12], p[8][11], r[36], c[36]);
HA HA_7(p[9][10], p[10][9], r[37], c[37]);
FA FA_30(p[0][20], p[1][19], p[2][18], r[38], c[38]);
FA FA_31(p[3][17], p[4][16], p[5][15], r[39], c[39]);
FA FA_32(p[6][14], p[7][13], p[8][12], r[40], c[40]);
FA FA_33(p[0][21], p[1][20], p[2][19], r[41], c[41]);
FA FA_34(p[3][18], p[4][17], p[5][16], r[42], c[42]);
FA FA_35(p[6][15], p[7][14], p[8][13], r[43], c[43]);
FA FA_36(p[0][22], p[1][21], p[2][20], r[44], c[44]);
FA FA_37(p[3][19], p[4][18], p[5][17], r[45], c[45]);
FA FA_38(p[6][16], p[7][15], p[8][14], r[46], c[46]);
HA HA_8(p[9][13], p[10][12], r[47], c[47]);
FA FA_39(p[0][23], p[1][22], p[2][21], r[48], c[48]);
FA FA_40(p[3][20], p[4][19], p[5][18], r[49], c[49]);
FA FA_41(p[6][17], p[7][16], p[8][15], r[50], c[50]);
FA FA_42(p[0][24], p[1][23], p[2][22], r[51], c[51]);
FA FA_43(p[3][21], p[4][20], p[5][19], r[52], c[52]);
FA FA_44(p[6][18], p[7][17], p[8][16], r[53], c[53]);
FA FA_45(p[0][25], p[1][24], p[2][23], r[54], c[54]);
FA FA_46(p[3][22], p[4][21], p[5][20], r[55], c[55]);
FA FA_47(p[6][19], p[7][18], p[8][17], r[56], c[56]);
HA HA_9(p[9][16], p[10][15], r[57], c[57]);
FA FA_48(p[0][26], p[1][25], p[2][24], r[58], c[58]);
FA FA_49(p[3][23], p[4][22], p[5][21], r[59], c[59]);
FA FA_50(p[6][20], p[7][19], p[8][18], r[60], c[60]);
FA FA_51(p[9][17], p[10][16], p[11][15], r[61], c[61]);
FA FA_52(p[0][27], p[1][26], p[2][25], r[62], c[62]);
FA FA_53(p[3][24], p[4][23], p[5][22], r[63], c[63]);
FA FA_54(p[6][21], p[7][20], p[8][19], r[64], c[64]);
FA FA_55(p[9][18], p[10][17], p[11][16], r[65], c[65]);
HA HA_10(p[12][15], p[13][14], r[66], c[66]);
FA FA_56(p[0][28], p[1][27], p[2][26], r[67], c[67]);
FA FA_57(p[3][25], p[4][24], p[5][23], r[68], c[68]);
FA FA_58(p[6][22], p[7][21], p[8][20], r[69], c[69]);
FA FA_59(p[9][19], p[10][18], p[11][17], r[70], c[70]);
FA FA_60(p[0][29], p[1][28], p[2][27], r[71], c[71]);
FA FA_61(p[3][26], p[4][25], p[5][24], r[72], c[72]);
FA FA_62(p[6][23], p[7][22], p[8][21], r[73], c[73]);
FA FA_63(p[9][20], p[10][19], p[11][18], r[74], c[74]);
FA FA_64(p[0][30], p[1][29], p[2][28], r[75], c[75]);
FA FA_65(p[3][27], p[4][26], p[5][25], r[76], c[76]);
FA FA_66(p[6][24], p[7][23], p[8][22], r[77], c[77]);
FA FA_67(p[9][21], p[10][20], p[11][19], r[78], c[78]);
HA HA_11(p[12][18], p[13][17], r[79], c[79]);
FA FA_68(p[0][31], p[1][30], p[2][29], r[80], c[80]);
FA FA_69(p[3][28], p[4][27], p[5][26], r[81], c[81]);
FA FA_70(p[6][25], p[7][24], p[8][23], r[82], c[82]);
FA FA_71(p[9][22], p[10][21], p[11][20], r[83], c[83]);
FA FA_72(p[1][31], p[2][30], p[3][29], r[84], c[84]);
FA FA_73(p[4][28], p[5][27], p[6][26], r[85], c[85]);
FA FA_74(p[7][25], p[8][24], p[9][23], r[86], c[86]);
FA FA_75(p[10][22], p[11][21], p[12][20], r[87], c[87]);
FA FA_76(p[2][31], p[3][30], p[4][29], r[88], c[88]);
FA FA_77(p[5][28], p[6][27], p[7][26], r[89], c[89]);
FA FA_78(p[8][25], p[9][24], p[10][23], r[90], c[90]);
FA FA_79(p[11][22], p[12][21], p[13][20], r[91], c[91]);
FA FA_80(p[3][31], p[4][30], p[5][29], r[92], c[92]);
FA FA_81(p[6][28], p[7][27], p[8][26], r[93], c[93]);
FA FA_82(p[9][25], p[10][24], p[11][23], r[94], c[94]);
FA FA_83(p[12][22], p[13][21], p[14][20], r[95], c[95]);
FA FA_84(p[4][31], p[5][30], p[6][29], r[96], c[96]);
FA FA_85(p[7][28], p[8][27], p[9][26], r[97], c[97]);
FA FA_86(p[10][25], p[11][24], p[12][23], r[98], c[98]);
FA FA_87(p[13][22], p[14][21], p[15][20], r[99], c[99]);
HA HA_12(p[16][19], p[17][18], r[100], c[100]);
FA FA_88(p[5][31], p[6][30], p[7][29], r[101], c[101]);
FA FA_89(p[8][28], p[9][27], p[10][26], r[102], c[102]);
FA FA_90(p[11][25], p[12][24], p[13][23], r[103], c[103]);
FA FA_91(p[14][22], p[15][21], p[16][20], r[104], c[104]);
HA HA_13(p[17][19], p[18][18], r[105], c[105]);
FA FA_92(p[6][31], p[7][30], p[8][29], r[106], c[106]);
FA FA_93(p[9][28], p[10][27], p[11][26], r[107], c[107]);
FA FA_94(p[12][25], p[13][24], p[14][23], r[108], c[108]);
FA FA_95(p[15][22], p[16][21], p[17][20], r[109], c[109]);
FA FA_96(p[7][31], p[8][30], p[9][29], r[110], c[110]);
FA FA_97(p[10][28], p[11][27], p[12][26], r[111], c[111]);
FA FA_98(p[13][25], p[14][24], p[15][23], r[112], c[112]);
HA HA_14(p[16][22], p[17][21], r[113], c[113]);
FA FA_99(p[8][31], p[9][30], p[10][29], r[114], c[114]);
FA FA_100(p[11][28], p[12][27], p[13][26], r[115], c[115]);
FA FA_101(p[14][25], p[15][24], p[16][23], r[116], c[116]);
FA FA_102(p[9][31], p[10][30], p[11][29], r[117], c[117]);
FA FA_103(p[12][28], p[13][27], p[14][26], r[118], c[118]);
FA FA_104(p[15][25], p[16][24], p[17][23], r[119], c[119]);
HA HA_15(p[18][22], p[19][21], r[120], c[120]);
FA FA_105(p[10][31], p[11][30], p[12][29], r[121], c[121]);
FA FA_106(p[13][28], p[14][27], p[15][26], r[122], c[122]);
FA FA_107(p[16][25], p[17][24], p[18][23], r[123], c[123]);
HA HA_16(p[19][22], p[20][21], r[124], c[124]);
FA FA_108(p[11][31], p[12][30], p[13][29], r[125], c[125]);
FA FA_109(p[14][28], p[15][27], p[16][26], r[126], c[126]);
FA FA_110(p[17][25], p[18][24], p[19][23], r[127], c[127]);
FA FA_111(p[12][31], p[13][30], p[14][29], r[128], c[128]);
FA FA_112(p[15][28], p[16][27], p[17][26], r[129], c[129]);
FA FA_113(p[18][25], p[19][24], p[20][23], r[130], c[130]);
HA HA_17(p[21][22], p[22][21], r[131], c[131]);
FA FA_114(p[13][31], p[14][30], p[15][29], r[132], c[132]);
FA FA_115(p[16][28], p[17][27], p[18][26], r[133], c[133]);
FA FA_116(p[19][25], p[20][24], p[21][23], r[134], c[134]);
HA HA_18(p[22][22], p[23][21], r[135], c[135]);
FA FA_117(p[14][31], p[15][30], p[16][29], r[136], c[136]);
FA FA_118(p[17][28], p[18][27], p[19][26], r[137], c[137]);
FA FA_119(p[20][25], p[21][24], p[22][23], r[138], c[138]);
FA FA_120(p[15][31], p[16][30], p[17][29], r[139], c[139]);
FA FA_121(p[18][28], p[19][27], p[20][26], r[140], c[140]);
HA HA_19(p[21][25], p[22][24], r[141], c[141]);
FA FA_122(p[16][31], p[17][30], p[18][29], r[142], c[142]);
FA FA_123(p[19][28], p[20][27], p[21][26], r[143], c[143]);
FA FA_124(p[17][31], p[18][30], p[19][29], r[144], c[144]);
FA FA_125(p[20][28], p[21][27], p[22][26], r[145], c[145]);
HA HA_20(p[23][25], p[24][24], r[146], c[146]);
FA FA_126(p[18][31], p[19][30], p[20][29], r[147], c[147]);
FA FA_127(p[21][28], p[22][27], p[23][26], r[148], c[148]);
HA HA_21(p[24][25], p[25][24], r[149], c[149]);
FA FA_128(p[19][31], p[20][30], p[21][29], r[150], c[150]);
FA FA_129(p[22][28], p[23][27], p[24][26], r[151], c[151]);
FA FA_130(p[20][31], p[21][30], p[22][29], r[152], c[152]);
FA FA_131(p[23][28], p[24][27], p[25][26], r[153], c[153]);
HA HA_22(p[26][25], p[27][24], r[154], c[154]);
FA FA_132(p[21][31], p[22][30], p[23][29], r[155], c[155]);
FA FA_133(p[24][28], p[25][27], p[26][26], r[156], c[156]);
HA HA_23(p[27][25], p[28][24], r[157], c[157]);
FA FA_134(p[22][31], p[23][30], p[24][29], r[158], c[158]);
FA FA_135(p[25][28], p[26][27], p[27][26], r[159], c[159]);
FA FA_136(p[23][31], p[24][30], p[25][29], r[160], c[160]);
HA HA_24(p[26][28], p[27][27], r[161], c[161]);
FA FA_137(p[24][31], p[25][30], p[26][29], r[162], c[162]);
FA FA_138(p[25][31], p[26][30], p[27][29], r[163], c[163]);
HA HA_25(p[28][28], p[29][27], r[164], c[164]);
FA FA_139(p[26][31], p[27][30], p[28][29], r[165], c[165]);
HA HA_26(p[29][28], p[30][27], r[166], c[166]);
FA FA_140(p[27][31], p[28][30], p[29][29], r[167], c[167]);
FA FA_141(p[28][31], p[29][30], p[30][29], r[168], c[168]);
HA HA_27(p[31][28], c[167], r[169], c[169]);
FA FA_142(p[29][31], p[30][30], p[31][29], r[170], c[170]);
HA HA_28(c[168], c[169], r[171], c[171]);
FA FA_143(p[30][31], p[31][30], c[170], r[172], c[172]);
HA HA_29(p[31][31], c[172], r[173], c[173]);
HA HA_30(1'b1, c[173], r[174], c[174]);
HA HA_31(c[0], r[1], r[175], c[175]);
FA FA_144(r[2], r[3], c[175], r[176], c[176]);
FA FA_145(p[3][1], p[4][0], c[2], r[177], c[177]);
FA FA_146(p[3][2], p[4][1], p[5][0], r[178], c[178]);
FA FA_147(p[5][1], p[6][0], c[5], r[179], c[179]);
FA FA_148(p[3][4], p[4][3], p[5][2], r[180], c[180]);
FA FA_149(p[3][5], p[4][4], p[5][3], r[181], c[181]);
FA FA_150(p[5][4], p[6][3], p[7][2], r[182], c[182]);
FA FA_151(p[6][4], p[7][3], p[8][2], r[183], c[183]);
FA FA_152(p[8][3], p[9][2], p[10][1], r[184], c[184]);
FA FA_153(p[6][6], p[7][5], p[8][4], r[185], c[185]);
FA FA_154(p[9][3], p[10][2], p[11][1], r[186], c[186]);
FA FA_155(p[6][7], p[7][6], p[8][5], r[187], c[187]);
FA FA_156(p[9][4], p[10][3], p[11][2], r[188], c[188]);
HA HA_32(p[12][1], p[13][0], r[189], c[189]);
FA FA_157(p[8][6], p[9][5], p[10][4], r[190], c[190]);
FA FA_158(p[11][3], p[12][2], p[13][1], r[191], c[191]);
FA FA_159(p[6][9], p[7][8], p[8][7], r[192], c[192]);
FA FA_160(p[9][6], p[10][5], p[11][4], r[193], c[193]);
HA HA_33(p[12][3], p[13][2], r[194], c[194]);
FA FA_161(p[6][10], p[7][9], p[8][8], r[195], c[195]);
FA FA_162(p[9][7], p[10][6], p[11][5], r[196], c[196]);
FA FA_163(p[8][9], p[9][8], p[10][7], r[197], c[197]);
FA FA_164(p[11][6], p[12][5], p[13][4], r[198], c[198]);
HA HA_34(p[14][3], p[15][2], r[199], c[199]);
FA FA_165(p[9][9], p[10][8], p[11][7], r[200], c[200]);
FA FA_166(p[12][6], p[13][5], p[14][4], r[201], c[201]);
FA FA_167(p[11][8], p[12][7], p[13][6], r[202], c[202]);
FA FA_168(p[14][5], p[15][4], p[16][3], r[203], c[203]);
FA FA_169(p[9][11], p[10][10], p[11][9], r[204], c[204]);
FA FA_170(p[12][8], p[13][7], p[14][6], r[205], c[205]);
FA FA_171(p[15][5], p[16][4], p[17][3], r[206], c[206]);
FA FA_172(p[9][12], p[10][11], p[11][10], r[207], c[207]);
FA FA_173(p[12][9], p[13][8], p[14][7], r[208], c[208]);
FA FA_174(p[15][6], p[16][5], p[17][4], r[209], c[209]);
FA FA_175(p[11][11], p[12][10], p[13][9], r[210], c[210]);
FA FA_176(p[14][8], p[15][7], p[16][6], r[211], c[211]);
FA FA_177(p[17][5], p[18][4], p[19][3], r[212], c[212]);
FA FA_178(p[9][14], p[10][13], p[11][12], r[213], c[213]);
FA FA_179(p[12][11], p[13][10], p[14][9], r[214], c[214]);
FA FA_180(p[15][8], p[16][7], p[17][6], r[215], c[215]);
FA FA_181(p[9][15], p[10][14], p[11][13], r[216], c[216]);
FA FA_182(p[12][12], p[13][11], p[14][10], r[217], c[217]);
FA FA_183(p[15][9], p[16][8], p[17][7], r[218], c[218]);
FA FA_184(p[11][14], p[12][13], p[13][12], r[219], c[219]);
FA FA_185(p[14][11], p[15][10], p[16][9], r[220], c[220]);
FA FA_186(p[17][8], p[18][7], p[19][6], r[221], c[221]);
FA FA_187(p[12][14], p[13][13], p[14][12], r[222], c[222]);
FA FA_188(p[15][11], p[16][10], p[17][9], r[223], c[223]);
FA FA_189(p[18][8], p[19][7], p[20][6], r[224], c[224]);
HA HA_35(p[21][5], p[22][4], r[225], c[225]);
FA FA_190(p[14][13], p[15][12], p[16][11], r[226], c[226]);
FA FA_191(p[17][10], p[18][9], p[19][8], r[227], c[227]);
FA FA_192(p[20][7], p[21][6], p[22][5], r[228], c[228]);
FA FA_193(p[12][16], p[13][15], p[14][14], r[229], c[229]);
FA FA_194(p[15][13], p[16][12], p[17][11], r[230], c[230]);
FA FA_195(p[18][10], p[19][9], p[20][8], r[231], c[231]);
HA HA_36(p[21][7], p[22][6], r[232], c[232]);
FA FA_196(p[12][17], p[13][16], p[14][15], r[233], c[233]);
FA FA_197(p[15][14], p[16][13], p[17][12], r[234], c[234]);
FA FA_198(p[18][11], p[19][10], p[20][9], r[235], c[235]);
FA FA_199(p[21][8], p[22][7], p[23][6], r[236], c[236]);
FA FA_200(p[14][16], p[15][15], p[16][14], r[237], c[237]);
FA FA_201(p[17][13], p[18][12], p[19][11], r[238], c[238]);
FA FA_202(p[20][10], p[21][9], p[22][8], r[239], c[239]);
FA FA_203(p[23][7], p[24][6], p[25][5], r[240], c[240]);
FA FA_204(p[12][19], p[13][18], p[14][17], r[241], c[241]);
FA FA_205(p[15][16], p[16][15], p[17][14], r[242], c[242]);
FA FA_206(p[18][13], p[19][12], p[20][11], r[243], c[243]);
FA FA_207(p[21][10], p[22][9], p[23][8], r[244], c[244]);
FA FA_208(p[13][19], p[14][18], p[15][17], r[245], c[245]);
FA FA_209(p[16][16], p[17][15], p[18][14], r[246], c[246]);
FA FA_210(p[19][13], p[20][12], p[21][11], r[247], c[247]);
FA FA_211(p[22][10], p[23][9], p[24][8], r[248], c[248]);
HA HA_37(p[25][7], p[26][6], r[249], c[249]);
FA FA_212(p[14][19], p[15][18], p[16][17], r[250], c[250]);
FA FA_213(p[17][16], p[18][15], p[19][14], r[251], c[251]);
FA FA_214(p[20][13], p[21][12], p[22][11], r[252], c[252]);
FA FA_215(p[23][10], p[24][9], p[25][8], r[253], c[253]);
FA FA_216(p[15][19], p[16][18], p[17][17], r[254], c[254]);
FA FA_217(p[18][16], p[19][15], p[20][14], r[255], c[255]);
FA FA_218(p[21][13], p[22][12], p[23][11], r[256], c[256]);
HA HA_38(p[24][10], p[25][9], r[257], c[257]);
FA FA_219(p[18][17], p[19][16], p[20][15], r[258], c[258]);
FA FA_220(p[21][14], p[22][13], p[23][12], r[259], c[259]);
FA FA_221(p[24][11], p[25][10], p[26][9], r[260], c[260]);
FA FA_222(p[19][17], p[20][16], p[21][15], r[261], c[261]);
FA FA_223(p[22][14], p[23][13], p[24][12], r[262], c[262]);
FA FA_224(p[25][11], p[26][10], p[27][9], r[263], c[263]);
HA HA_39(p[28][8], p[29][7], r[264], c[264]);
FA FA_225(p[18][19], p[19][18], p[20][17], r[265], c[265]);
FA FA_226(p[21][16], p[22][15], p[23][14], r[266], c[266]);
FA FA_227(p[24][13], p[25][12], p[26][11], r[267], c[267]);
FA FA_228(p[18][20], p[19][19], p[20][18], r[268], c[268]);
FA FA_229(p[21][17], p[22][16], p[23][15], r[269], c[269]);
FA FA_230(p[24][14], p[25][13], p[26][12], r[270], c[270]);
FA FA_231(p[17][22], p[18][21], p[19][20], r[271], c[271]);
FA FA_232(p[20][19], p[21][18], p[22][17], r[272], c[272]);
FA FA_233(p[23][16], p[24][15], p[25][14], r[273], c[273]);
FA FA_234(p[20][20], p[21][19], p[22][18], r[274], c[274]);
FA FA_235(p[23][17], p[24][16], p[25][15], r[275], c[275]);
FA FA_236(p[26][14], p[27][13], p[28][12], r[276], c[276]);
FA FA_237(p[21][20], p[22][19], p[23][18], r[277], c[277]);
FA FA_238(p[24][17], p[25][16], p[26][15], r[278], c[278]);
FA FA_239(p[27][14], p[28][13], p[29][12], r[279], c[279]);
FA FA_240(p[20][22], p[21][21], p[22][20], r[280], c[280]);
FA FA_241(p[23][19], p[24][18], p[25][17], r[281], c[281]);
FA FA_242(p[26][16], p[27][15], p[28][14], r[282], c[282]);
FA FA_243(p[23][20], p[24][19], p[25][18], r[283], c[283]);
FA FA_244(p[26][17], p[27][16], p[28][15], r[284], c[284]);
FA FA_245(p[24][20], p[25][19], p[26][18], r[285], c[285]);
FA FA_246(p[27][17], p[28][16], p[29][15], r[286], c[286]);
FA FA_247(p[23][22], p[24][21], p[25][20], r[287], c[287]);
FA FA_248(p[26][19], p[27][18], p[28][17], r[288], c[288]);
FA FA_249(p[23][23], p[24][22], p[25][21], r[289], c[289]);
FA FA_250(p[26][20], p[27][19], p[28][18], r[290], c[290]);
HA HA_40(p[29][17], p[30][16], r[291], c[291]);
FA FA_251(p[22][25], p[23][24], p[24][23], r[292], c[292]);
FA FA_252(p[25][22], p[26][21], p[27][20], r[293], c[293]);
FA FA_253(p[25][23], p[26][22], p[27][21], r[294], c[294]);
FA FA_254(p[28][20], p[29][19], p[30][18], r[295], c[295]);
HA HA_41(p[31][17], c[142], r[296], c[296]);
FA FA_255(p[26][23], p[27][22], p[28][21], r[297], c[297]);
FA FA_256(p[29][20], p[30][19], p[31][18], r[298], c[298]);
FA FA_257(p[25][25], p[26][24], p[27][23], r[299], c[299]);
FA FA_258(p[28][22], p[29][21], p[30][20], r[300], c[300]);
HA HA_42(p[31][19], c[147], r[301], c[301]);
FA FA_259(p[28][23], p[29][22], p[30][21], r[302], c[302]);
FA FA_260(p[31][20], c[150], c[151], r[303], c[303]);
FA FA_261(p[29][23], p[30][22], p[31][21], r[304], c[304]);
HA HA_43(c[152], c[153], r[305], c[305]);
FA FA_262(p[28][25], p[29][24], p[30][23], r[306], c[306]);
HA HA_44(p[31][22], c[155], r[307], c[307]);
FA FA_263(p[28][26], p[29][25], p[30][24], r[308], c[308]);
FA FA_264(p[27][28], p[28][27], p[29][26], r[309], c[309]);
FA FA_265(p[30][26], p[31][25], c[162], r[310], c[310]);
FA FA_266(p[31][26], c[163], c[164], r[311], c[311]);
FA FA_267(p[30][28], p[31][27], c[165], r[312], c[312]);
FA FA_268(r[168], r[169], c[312], r[313], c[313]);
FA FA_269(r[170], r[171], c[313], r[314], c[314]);
FA FA_270(c[171], r[172], c[314], r[315], c[315]);
HA HA_45(r[173], c[315], r[316], c[316]);
HA HA_46(r[174], c[316], r[317], c[317]);
FA FA_271(c[3], r[4], c[176], r[318], c[318]);
FA FA_272(c[4], r[5], c[177], r[319], c[319]);
HA HA_47(r[178], c[318], r[320], c[320]);
FA FA_273(r[6], r[7], c[178], r[321], c[321]);
FA FA_274(p[6][1], p[7][0], c[6], r[322], c[322]);
HA HA_48(c[7], r[8], r[323], c[323]);
FA FA_275(p[6][2], p[7][1], p[8][0], r[324], c[324]);
FA FA_276(p[8][1], p[9][0], c[9], r[325], c[325]);
HA HA_49(r[10], r[11], r[326], c[326]);
FA FA_277(p[9][1], p[10][0], c[10], r[327], c[327]);
FA FA_278(p[11][0], c[12], c[13], r[328], c[328]);
FA FA_279(p[12][0], c[14], c[15], r[329], c[329]);
FA FA_280(c[17], c[18], r[19], r[330], c[330]);
FA FA_281(p[14][0], c[19], c[20], r[331], c[331]);
FA FA_282(r[21], r[22], r[23], r[332], c[332]);
FA FA_283(p[14][1], p[15][0], c[21], r[333], c[333]);
FA FA_284(c[22], c[23], r[24], r[334], c[334]);
HA HA_50(r[25], c[190], r[335], c[335]);
FA FA_285(p[12][4], p[13][3], p[14][2], r[336], c[336]);
FA FA_286(p[15][1], p[16][0], c[24], r[337], c[337]);
HA HA_51(c[25], r[26], r[338], c[338]);
FA FA_287(p[16][1], p[17][0], c[26], r[339], c[339]);
FA FA_288(c[27], r[28], r[29], r[340], c[340]);
FA FA_289(p[15][3], p[16][2], p[17][1], r[341], c[341]);
FA FA_290(p[18][0], c[28], c[29], r[342], c[342]);
HA HA_52(c[30], r[31], r[343], c[343]);
FA FA_291(p[17][2], p[18][1], p[19][0], r[344], c[344]);
FA FA_292(c[31], c[32], c[33], r[345], c[345]);
HA HA_53(r[34], r[35], r[346], c[346]);
FA FA_293(p[18][2], p[19][1], p[20][0], r[347], c[347]);
FA FA_294(c[34], c[35], c[36], r[348], c[348]);
FA FA_295(p[18][3], p[19][2], p[20][1], r[349], c[349]);
FA FA_296(p[21][0], c[38], c[39], r[350], c[350]);
FA FA_297(p[20][2], p[21][1], p[22][0], r[351], c[351]);
FA FA_298(c[41], c[42], c[43], r[352], c[352]);
FA FA_299(p[18][5], p[19][4], p[20][3], r[353], c[353]);
FA FA_300(p[21][2], p[22][1], p[23][0], r[354], c[354]);
FA FA_301(c[44], c[45], c[46], r[355], c[355]);
FA FA_302(p[18][6], p[19][5], p[20][4], r[356], c[356]);
FA FA_303(p[21][3], p[22][2], p[23][1], r[357], c[357]);
FA FA_304(p[24][0], c[48], c[49], r[358], c[358]);
FA FA_305(p[20][5], p[21][4], p[22][3], r[359], c[359]);
FA FA_306(p[23][2], p[24][1], p[25][0], r[360], c[360]);
FA FA_307(c[51], c[52], c[53], r[361], c[361]);
FA FA_308(p[23][3], p[24][2], p[25][1], r[362], c[362]);
FA FA_309(p[26][0], c[54], c[55], r[363], c[363]);
FA FA_310(c[56], c[57], r[58], r[364], c[364]);
FA FA_311(p[23][4], p[24][3], p[25][2], r[365], c[365]);
FA FA_312(p[26][1], p[27][0], c[58], r[366], c[366]);
FA FA_313(c[59], c[60], c[61], r[367], c[367]);
FA FA_314(p[23][5], p[24][4], p[25][3], r[368], c[368]);
FA FA_315(p[26][2], p[27][1], p[28][0], r[369], c[369]);
FA FA_316(c[62], c[63], c[64], r[370], c[370]);
FA FA_317(p[24][5], p[25][4], p[26][3], r[371], c[371]);
FA FA_318(p[27][2], p[28][1], p[29][0], r[372], c[372]);
FA FA_319(c[67], c[68], c[69], r[373], c[373]);
FA FA_320(p[26][4], p[27][3], p[28][2], r[374], c[374]);
FA FA_321(p[29][1], p[30][0], c[71], r[375], c[375]);
FA FA_322(c[72], c[73], c[74], r[376], c[376]);
FA FA_323(p[24][7], p[25][6], p[26][5], r[377], c[377]);
FA FA_324(p[27][4], p[28][3], p[29][2], r[378], c[378]);
FA FA_325(p[30][1], p[31][0], c[75], r[379], c[379]);
FA FA_326(p[27][5], p[28][4], p[29][3], r[380], c[380]);
FA FA_327(p[30][2], p[31][1], 1'b1, r[381], c[381]);
FA FA_328(c[80], c[81], c[82], r[382], c[382]);
HA HA_54(c[83], r[84], r[383], c[383]);
FA FA_329(p[26][7], p[27][6], p[28][5], r[384], c[384]);
FA FA_330(p[29][4], p[30][3], p[31][2], r[385], c[385]);
FA FA_331(c[84], c[85], c[86], r[386], c[386]);
FA FA_332(p[26][8], p[27][7], p[28][6], r[387], c[387]);
FA FA_333(p[29][5], p[30][4], p[31][3], r[388], c[388]);
FA FA_334(c[88], c[89], c[90], r[389], c[389]);
FA FA_335(p[27][8], p[28][7], p[29][6], r[390], c[390]);
FA FA_336(p[30][5], p[31][4], c[92], r[391], c[391]);
FA FA_337(c[93], c[94], c[95], r[392], c[392]);
FA FA_338(p[30][6], p[31][5], c[96], r[393], c[393]);
FA FA_339(c[97], c[98], c[99], r[394], c[394]);
FA FA_340(c[100], r[101], r[102], r[395], c[395]);
FA FA_341(p[27][10], p[28][9], p[29][8], r[396], c[396]);
FA FA_342(p[30][7], p[31][6], c[101], r[397], c[397]);
FA FA_343(c[102], c[103], c[104], r[398], c[398]);
FA FA_344(p[27][11], p[28][10], p[29][9], r[399], c[399]);
FA FA_345(p[30][8], p[31][7], c[106], r[400], c[400]);
FA FA_346(c[107], c[108], c[109], r[401], c[401]);
FA FA_347(p[26][13], p[27][12], p[28][11], r[402], c[402]);
FA FA_348(p[29][10], p[30][9], p[31][8], r[403], c[403]);
FA FA_349(c[110], c[111], c[112], r[404], c[404]);
FA FA_350(p[29][11], p[30][10], p[31][9], r[405], c[405]);
FA FA_351(c[114], c[115], c[116], r[406], c[406]);
FA FA_352(p[30][11], p[31][10], c[117], r[407], c[407]);
FA FA_353(c[118], c[119], c[120], r[408], c[408]);
FA FA_354(p[29][13], p[30][12], p[31][11], r[409], c[409]);
FA FA_355(c[121], c[122], c[123], r[410], c[410]);
FA FA_356(p[29][14], p[30][13], p[31][12], r[411], c[411]);
FA FA_357(c[125], c[126], c[127], r[412], c[412]);
HA HA_55(r[128], r[129], r[413], c[413]);
FA FA_358(p[30][14], p[31][13], c[128], r[414], c[414]);
FA FA_359(c[129], c[130], c[131], r[415], c[415]);
HA HA_56(r[132], r[133], r[416], c[416]);
FA FA_360(p[29][16], p[30][15], p[31][14], r[417], c[417]);
FA FA_361(c[132], c[133], c[134], r[418], c[418]);
HA HA_57(c[135], r[136], r[419], c[419]);
FA FA_362(p[31][15], c[136], c[137], r[420], c[420]);
FA FA_363(c[138], r[139], r[140], r[421], c[421]);
FA FA_364(p[28][19], p[29][18], p[30][17], r[422], c[422]);
FA FA_365(p[31][16], c[139], c[140], r[423], c[423]);
FA FA_366(c[143], r[144], r[145], r[424], c[424]);
HA HA_58(r[146], c[292], r[425], c[425]);
FA FA_367(c[144], c[145], c[146], r[426], c[426]);
FA FA_368(r[147], r[148], r[149], r[427], c[427]);
FA FA_369(c[148], c[149], r[150], r[428], c[428]);
HA HA_59(r[151], c[297], r[429], c[429]);
FA FA_370(r[152], r[153], r[154], r[430], c[430]);
FA FA_371(c[154], r[155], r[156], r[431], c[431]);
FA FA_372(c[156], c[157], r[158], r[432], c[432]);
FA FA_373(p[31][23], c[158], c[159], r[433], c[433]);
FA FA_374(p[30][25], p[31][24], c[160], r[434], c[434]);
HA HA_60(c[161], r[162], r[435], c[435]);
FA FA_375(r[163], r[164], c[309], r[436], c[436]);
FA FA_376(r[165], r[166], c[310], r[437], c[437]);
HA HA_61(r[311], c[436], r[438], c[438]);
FA FA_377(c[166], r[167], c[311], r[439], c[439]);
HA HA_62(r[313], c[439], r[440], c[440]);
HA HA_63(r[314], c[440], r[441], c[441]);
HA HA_64(r[315], c[441], r[442], c[442]);
HA HA_65(r[316], c[442], r[443], c[443]);
HA HA_66(r[317], c[443], r[444], c[444]);
HA HA_67(r[177], r[318], r[445], c[445]);
FA FA_378(r[319], r[320], c[445], r[446], c[446]);
FA FA_379(r[179], c[319], c[320], r[447], c[447]);
HA HA_68(r[321], c[446], r[448], c[448]);
FA FA_380(c[179], r[180], c[321], r[449], c[449]);
FA FA_381(c[8], r[9], c[180], r[450], c[450]);
HA HA_69(r[181], c[322], r[451], c[451]);
FA FA_382(c[181], r[182], c[324], r[452], c[452]);
FA FA_383(c[11], r[12], r[13], r[453], c[453]);
FA FA_384(r[14], r[15], r[16], r[454], c[454]);
HA HA_70(c[183], r[184], r[455], c[455]);
FA FA_385(c[16], r[17], r[18], r[456], c[456]);
FA FA_386(r[20], c[185], c[186], r[457], c[457]);
FA FA_387(c[187], c[188], c[189], r[458], c[458]);
FA FA_388(c[191], r[192], r[193], r[459], c[459]);
FA FA_389(r[27], c[192], c[193], r[460], c[460]);
FA FA_390(c[194], r[195], r[196], r[461], c[461]);
FA FA_391(r[30], c[195], c[196], r[462], c[462]);
FA FA_392(r[197], r[198], r[199], r[463], c[463]);
FA FA_393(r[32], r[33], c[197], r[464], c[464]);
FA FA_394(c[198], c[199], r[200], r[465], c[465]);
HA HA_71(r[201], c[339], r[466], c[466]);
FA FA_395(r[36], r[37], c[200], r[467], c[467]);
FA FA_396(c[201], r[202], r[203], r[468], c[468]);
FA FA_397(c[37], r[38], r[39], r[469], c[469]);
FA FA_398(r[40], c[202], c[203], r[470], c[470]);
FA FA_399(c[40], r[41], r[42], r[471], c[471]);
FA FA_400(r[43], c[204], c[205], r[472], c[472]);
FA FA_401(r[44], r[45], r[46], r[473], c[473]);
FA FA_402(r[47], c[207], c[208], r[474], c[474]);
FA FA_403(c[47], r[48], r[49], r[475], c[475]);
FA FA_404(r[50], c[210], c[211], r[476], c[476]);
HA HA_72(c[212], r[213], r[477], c[477]);
FA FA_405(c[50], r[51], r[52], r[478], c[478]);
FA FA_406(r[53], c[213], c[214], r[479], c[479]);
FA FA_407(r[54], r[55], r[56], r[480], c[480]);
FA FA_408(r[57], c[216], c[217], r[481], c[481]);
FA FA_409(r[59], r[60], r[61], r[482], c[482]);
FA FA_410(c[219], c[220], c[221], r[483], c[483]);
FA FA_411(r[62], r[63], r[64], r[484], c[484]);
FA FA_412(r[65], r[66], c[222], r[485], c[485]);
HA HA_73(c[223], c[224], r[486], c[486]);
FA FA_413(c[65], c[66], r[67], r[487], c[487]);
FA FA_414(r[68], r[69], r[70], r[488], c[488]);
FA FA_415(c[226], c[227], c[228], r[489], c[489]);
FA FA_416(c[70], r[71], r[72], r[490], c[490]);
FA FA_417(r[73], r[74], c[229], r[491], c[491]);
FA FA_418(c[230], c[231], c[232], r[492], c[492]);
FA FA_419(r[75], r[76], r[77], r[493], c[493]);
FA FA_420(r[78], r[79], c[233], r[494], c[494]);
FA FA_421(c[234], c[235], c[236], r[495], c[495]);
FA FA_422(c[76], c[77], c[78], r[496], c[496]);
FA FA_423(c[79], r[80], r[81], r[497], c[497]);
FA FA_424(r[82], r[83], c[237], r[498], c[498]);
FA FA_425(r[85], r[86], r[87], r[499], c[499]);
FA FA_426(c[241], c[242], c[243], r[500], c[500]);
FA FA_427(c[244], r[245], r[246], r[501], c[501]);
FA FA_428(c[87], r[88], r[89], r[502], c[502]);
FA FA_429(r[90], r[91], c[245], r[503], c[503]);
FA FA_430(c[246], c[247], c[248], r[504], c[504]);
FA FA_431(c[91], r[92], r[93], r[505], c[505]);
FA FA_432(r[94], r[95], c[250], r[506], c[506]);
FA FA_433(c[251], c[252], c[253], r[507], c[507]);
FA FA_434(r[96], r[97], r[98], r[508], c[508]);
FA FA_435(r[99], r[100], c[254], r[509], c[509]);
FA FA_436(c[255], c[256], c[257], r[510], c[510]);
FA FA_437(r[103], r[104], r[105], r[511], c[511]);
FA FA_438(c[258], c[259], c[260], r[512], c[512]);
FA FA_439(c[105], r[106], r[107], r[513], c[513]);
FA FA_440(r[108], r[109], c[261], r[514], c[514]);
HA HA_74(c[262], c[263], r[515], c[515]);
FA FA_441(r[110], r[111], r[112], r[516], c[516]);
FA FA_442(r[113], c[265], c[266], r[517], c[517]);
FA FA_443(c[113], r[114], r[115], r[518], c[518]);
FA FA_444(r[116], c[268], c[269], r[519], c[519]);
FA FA_445(r[117], r[118], r[119], r[520], c[520]);
FA FA_446(r[120], c[271], c[272], r[521], c[521]);
HA HA_75(c[273], r[274], r[522], c[522]);
FA FA_447(r[121], r[122], r[123], r[523], c[523]);
FA FA_448(r[124], c[274], c[275], r[524], c[524]);
HA HA_76(c[276], r[277], r[525], c[525]);
FA FA_449(c[124], r[125], r[126], r[526], c[526]);
FA FA_450(r[127], c[277], c[278], r[527], c[527]);
HA HA_77(c[279], r[280], r[528], c[528]);
FA FA_451(r[130], r[131], c[280], r[529], c[529]);
FA FA_452(c[281], c[282], r[283], r[530], c[530]);
FA FA_453(r[134], r[135], c[283], r[531], c[531]);
FA FA_454(c[284], r[285], r[286], r[532], c[532]);
HA HA_78(c[411], c[412], r[533], c[533]);
FA FA_455(r[137], r[138], c[285], r[534], c[534]);
FA FA_456(c[286], r[287], r[288], r[535], c[535]);
FA FA_457(r[141], c[287], c[288], r[536], c[536]);
FA FA_458(r[289], r[290], r[291], r[537], c[537]);
FA FA_459(c[141], r[142], r[143], r[538], c[538]);
FA FA_460(c[289], c[290], c[291], r[539], c[539]);
HA HA_79(r[292], r[293], r[540], c[540]);
FA FA_461(c[293], r[294], r[295], r[541], c[541]);
HA HA_80(r[296], c[422], r[542], c[542]);
FA FA_462(c[294], c[295], c[296], r[543], c[543]);
HA HA_81(r[297], r[298], r[544], c[544]);
FA FA_463(c[298], r[299], r[300], r[545], c[545]);
FA FA_464(c[299], c[300], c[301], r[546], c[546]);
FA FA_465(r[157], c[302], c[303], r[547], c[547]);
HA HA_82(r[304], r[305], r[548], c[548]);
FA FA_466(r[159], c[304], c[305], r[549], c[549]);
FA FA_467(r[160], r[161], c[306], r[550], c[550]);
HA HA_83(c[307], r[308], r[551], c[551]);
FA FA_468(c[308], r[309], c[433], r[552], c[552]);
FA FA_469(r[310], c[434], c[435], r[553], c[553]);
HA HA_84(r[436], c[552], r[554], c[554]);
FA FA_470(r[437], r[438], c[553], r[555], c[555]);
FA FA_471(r[312], c[437], c[438], r[556], c[556]);
HA HA_85(r[439], c[555], r[557], c[557]);
FA FA_472(r[440], c[556], c[557], r[558], c[558]);
HA HA_86(r[441], c[558], r[559], c[559]);
HA HA_87(r[442], c[559], r[560], c[560]);
HA HA_88(r[443], c[560], r[561], c[561]);
HA HA_89(r[444], c[561], r[562], c[562]);
HA HA_90(r[447], r[448], r[563], c[563]);
FA FA_473(r[322], r[323], c[447], r[564], c[564]);
FA FA_474(c[323], r[324], c[449], r[565], c[565]);
FA FA_475(r[325], r[326], c[450], r[566], c[566]);
FA FA_476(c[182], r[183], c[325], r[567], c[567]);
HA HA_91(c[326], r[327], r[568], c[568]);
FA FA_477(c[327], r[328], c[453], r[569], c[569]);
FA FA_478(c[184], r[185], r[186], r[570], c[570]);
FA FA_479(r[187], r[188], r[189], r[571], c[571]);
HA HA_92(c[329], r[330], r[572], c[572]);
FA FA_480(r[190], r[191], c[330], r[573], c[573]);
FA FA_481(r[194], c[331], c[332], r[574], c[574]);
FA FA_482(c[333], c[334], c[335], r[575], c[575]);
FA FA_483(c[336], c[337], c[338], r[576], c[576]);
FA FA_484(c[340], r[341], r[342], r[577], c[577]);
FA FA_485(c[341], c[342], c[343], r[578], c[578]);
FA FA_486(r[344], r[345], r[346], r[579], c[579]);
FA FA_487(r[204], r[205], r[206], r[580], c[580]);
FA FA_488(c[344], c[345], c[346], r[581], c[581]);
HA HA_93(r[347], r[348], r[582], c[582]);
FA FA_489(c[206], r[207], r[208], r[583], c[583]);
FA FA_490(r[209], c[347], c[348], r[584], c[584]);
FA FA_491(c[209], r[210], r[211], r[585], c[585]);
FA FA_492(r[212], c[349], c[350], r[586], c[586]);
HA HA_94(r[351], r[352], r[587], c[587]);
FA FA_493(r[214], r[215], c[351], r[588], c[588]);
FA FA_494(c[352], r[353], r[354], r[589], c[589]);
FA FA_495(c[215], r[216], r[217], r[590], c[590]);
FA FA_496(r[218], c[353], c[354], r[591], c[591]);
HA HA_95(c[355], r[356], r[592], c[592]);
FA FA_497(c[218], r[219], r[220], r[593], c[593]);
FA FA_498(r[221], c[356], c[357], r[594], c[594]);
HA HA_96(c[358], r[359], r[595], c[595]);
FA FA_499(r[222], r[223], r[224], r[596], c[596]);
FA FA_500(r[225], c[359], c[360], r[597], c[597]);
HA HA_97(c[361], r[362], r[598], c[598]);
FA FA_501(c[225], r[226], r[227], r[599], c[599]);
FA FA_502(r[228], c[362], c[363], r[600], c[600]);
FA FA_503(r[229], r[230], r[231], r[601], c[601]);
FA FA_504(r[232], c[365], c[366], r[602], c[602]);
FA FA_505(r[233], r[234], r[235], r[603], c[603]);
FA FA_506(r[236], c[368], c[369], r[604], c[604]);
FA FA_507(r[237], r[238], r[239], r[605], c[605]);
FA FA_508(r[240], c[371], c[372], r[606], c[606]);
FA FA_509(c[238], c[239], c[240], r[607], c[607]);
FA FA_510(r[241], r[242], r[243], r[608], c[608]);
FA FA_511(r[244], c[374], c[375], r[609], c[609]);
FA FA_512(r[247], r[248], r[249], r[610], c[610]);
FA FA_513(c[377], c[378], c[379], r[611], c[611]);
FA FA_514(c[249], r[250], r[251], r[612], c[612]);
FA FA_515(r[252], r[253], c[380], r[613], c[613]);
HA HA_98(c[381], c[382], r[614], c[614]);
FA FA_516(r[254], r[255], r[256], r[615], c[615]);
FA FA_517(r[257], c[384], c[385], r[616], c[616]);
FA FA_518(r[258], r[259], r[260], r[617], c[617]);
FA FA_519(c[387], c[388], c[389], r[618], c[618]);
HA HA_99(r[390], r[391], r[619], c[619]);
FA FA_520(r[261], r[262], r[263], r[620], c[620]);
FA FA_521(r[264], c[390], c[391], r[621], c[621]);
FA FA_522(c[264], r[265], r[266], r[622], c[622]);
FA FA_523(r[267], c[393], c[394], r[623], c[623]);
HA HA_100(c[395], r[396], r[624], c[624]);
FA FA_524(c[267], r[268], r[269], r[625], c[625]);
FA FA_525(r[270], c[396], c[397], r[626], c[626]);
FA FA_526(c[270], r[271], r[272], r[627], c[627]);
FA FA_527(r[273], c[399], c[400], r[628], c[628]);
FA FA_528(r[275], r[276], c[402], r[629], c[629]);
FA FA_529(c[403], c[404], r[405], r[630], c[630]);
HA HA_101(r[406], c[518], r[631], c[631]);
FA FA_530(r[278], r[279], c[405], r[632], c[632]);
FA FA_531(c[406], r[407], r[408], r[633], c[633]);
FA FA_532(r[281], r[282], c[407], r[634], c[634]);
FA FA_533(c[408], r[409], r[410], r[635], c[635]);
HA HA_102(c[523], c[524], r[636], c[636]);
FA FA_534(r[284], c[409], c[410], r[637], c[637]);
FA FA_535(r[411], r[412], r[413], r[638], c[638]);
HA HA_103(c[526], c[527], r[639], c[639]);
FA FA_536(c[413], r[414], r[415], r[640], c[640]);
FA FA_537(r[416], c[529], c[530], r[641], c[641]);
FA FA_538(c[414], c[415], c[416], r[642], c[642]);
FA FA_539(r[417], r[418], r[419], r[643], c[643]);
FA FA_540(c[417], c[418], c[419], r[644], c[644]);
HA HA_104(r[420], r[421], r[645], c[645]);
FA FA_541(c[420], c[421], r[422], r[646], c[646]);
HA HA_105(r[423], c[536], r[647], c[647]);
FA FA_542(c[423], r[424], r[425], r[648], c[648]);
FA FA_543(c[424], c[425], r[426], r[649], c[649]);
FA FA_544(r[301], c[426], c[427], r[650], c[650]);
FA FA_545(r[302], r[303], c[428], r[651], c[651]);
HA HA_106(c[429], r[430], r[652], c[652]);
FA FA_546(c[430], r[431], c[546], r[653], c[653]);
FA FA_547(r[306], r[307], c[431], r[654], c[654]);
HA HA_107(r[432], c[547], r[655], c[655]);
FA FA_548(c[432], r[433], c[549], r[656], c[656]);
FA FA_549(r[434], r[435], c[550], r[657], c[657]);
FA FA_550(r[553], r[554], c[657], r[658], c[658]);
FA FA_551(c[554], r[555], c[658], r[659], c[659]);
FA FA_552(r[556], r[557], c[659], r[660], c[660]);
HA HA_108(r[558], c[660], r[661], c[661]);
HA HA_109(r[559], c[661], r[662], c[662]);
HA HA_110(r[560], c[662], r[663], c[663]);
HA HA_111(r[561], c[663], r[664], c[664]);
HA HA_112(r[562], c[664], r[665], c[665]);
FA FA_553(c[448], r[449], c[563], r[666], c[666]);
FA FA_554(r[450], r[451], c[564], r[667], c[667]);
HA HA_113(r[565], c[666], r[668], c[668]);
FA FA_555(c[451], r[452], c[565], r[669], c[669]);
FA FA_556(c[452], r[453], c[566], r[670], c[670]);
FA FA_557(r[454], r[455], c[567], r[671], c[671]);
FA FA_558(c[328], r[329], c[454], r[672], c[672]);
HA HA_114(c[455], r[456], r[673], c[673]);
FA FA_559(c[456], r[457], c[570], r[674], c[674]);
FA FA_560(r[331], r[332], c[457], r[675], c[675]);
HA HA_115(r[458], c[571], r[676], c[676]);
FA FA_561(r[333], r[334], r[335], r[677], c[677]);
FA FA_562(r[336], r[337], r[338], r[678], c[678]);
FA FA_563(r[339], r[340], c[460], r[679], c[679]);
FA FA_564(r[343], c[462], c[463], r[680], c[680]);
FA FA_565(c[464], c[465], c[466], r[681], c[681]);
FA FA_566(c[467], c[468], r[469], r[682], c[682]);
FA FA_567(r[349], r[350], c[469], r[683], c[683]);
FA FA_568(c[470], r[471], r[472], r[684], c[684]);
FA FA_569(c[471], c[472], r[473], r[685], c[685]);
HA HA_116(r[474], c[583], r[686], c[686]);
FA FA_570(r[355], c[473], c[474], r[687], c[687]);
FA FA_571(r[475], r[476], r[477], r[688], c[688]);
FA FA_572(r[357], r[358], c[475], r[689], c[689]);
FA FA_573(c[476], c[477], r[478], r[690], c[690]);
HA HA_117(r[479], c[588], r[691], c[691]);
FA FA_574(r[360], r[361], c[478], r[692], c[692]);
FA FA_575(c[479], r[480], r[481], r[693], c[693]);
FA FA_576(r[363], r[364], c[480], r[694], c[694]);
FA FA_577(c[481], r[482], r[483], r[695], c[695]);
HA HA_118(c[593], c[594], r[696], c[696]);
FA FA_578(c[364], r[365], r[366], r[697], c[697]);
FA FA_579(r[367], c[482], c[483], r[698], c[698]);
HA HA_119(r[484], r[485], r[699], c[699]);
FA FA_580(c[367], r[368], r[369], r[700], c[700]);
FA FA_581(r[370], c[484], c[485], r[701], c[701]);
HA HA_120(c[486], r[487], r[702], c[702]);
FA FA_582(c[370], r[371], r[372], r[703], c[703]);
FA FA_583(r[373], c[487], c[488], r[704], c[704]);
HA HA_121(c[489], r[490], r[705], c[705]);
FA FA_584(c[373], r[374], r[375], r[706], c[706]);
FA FA_585(r[376], c[490], c[491], r[707], c[707]);
HA HA_122(c[492], r[493], r[708], c[708]);
FA FA_586(c[376], r[377], r[378], r[709], c[709]);
FA FA_587(r[379], c[493], c[494], r[710], c[710]);
FA FA_588(r[380], r[381], r[382], r[711], c[711]);
FA FA_589(r[383], c[496], c[497], r[712], c[712]);
HA HA_123(c[498], r[499], r[713], c[713]);
FA FA_590(c[383], r[384], r[385], r[714], c[714]);
FA FA_591(r[386], c[499], c[500], r[715], c[715]);
FA FA_592(c[386], r[387], r[388], r[716], c[716]);
FA FA_593(r[389], c[502], c[503], r[717], c[717]);
HA HA_124(c[504], r[505], r[718], c[718]);
FA FA_594(r[392], c[505], c[506], r[719], c[719]);
FA FA_595(c[507], r[508], r[509], r[720], c[720]);
FA FA_596(c[392], r[393], r[394], r[721], c[721]);
FA FA_597(r[395], c[508], c[509], r[722], c[722]);
FA FA_598(r[397], r[398], c[511], r[723], c[723]);
FA FA_599(c[512], r[513], r[514], r[724], c[724]);
HA HA_125(r[515], c[620], r[725], c[725]);
FA FA_600(c[398], r[399], r[400], r[726], c[726]);
FA FA_601(r[401], c[513], c[514], r[727], c[727]);
HA HA_126(c[515], r[516], r[728], c[728]);
FA FA_602(c[401], r[402], r[403], r[729], c[729]);
FA FA_603(r[404], c[516], c[517], r[730], c[730]);
FA FA_604(c[519], r[520], r[521], r[731], c[731]);
HA HA_127(r[522], c[627], r[732], c[732]);
FA FA_605(c[520], c[521], c[522], r[733], c[733]);
FA FA_606(r[523], r[524], r[525], r[734], c[734]);
FA FA_607(c[525], r[526], r[527], r[735], c[735]);
HA HA_128(r[528], c[632], r[736], c[736]);
FA FA_608(c[528], r[529], r[530], r[737], c[737]);
HA HA_129(c[634], c[635], r[738], c[738]);
FA FA_609(r[531], r[532], r[533], r[739], c[739]);
FA FA_610(c[531], c[532], c[533], r[740], c[740]);
FA FA_611(c[534], c[535], r[536], r[741], c[741]);
FA FA_612(c[537], r[538], r[539], r[742], c[742]);
FA FA_613(c[538], c[539], c[540], r[743], c[743]);
FA FA_614(r[427], c[541], c[542], r[744], c[744]);
HA HA_130(r[543], r[544], r[745], c[745]);
FA FA_615(r[428], r[429], c[543], r[746], c[746]);
FA FA_616(c[545], r[546], c[650], r[747], c[747]);
FA FA_617(r[547], r[548], c[651], r[748], c[748]);
FA FA_618(c[548], r[549], c[653], r[749], c[749]);
FA FA_619(r[550], r[551], c[654], r[750], c[750]);
FA FA_620(c[551], r[552], c[656], r[751], c[751]);
HA HA_131(r[657], c[750], r[752], c[752]);
FA FA_621(r[658], c[751], c[752], r[753], c[753]);
HA HA_132(r[659], c[753], r[754], c[754]);
HA HA_133(r[660], c[754], r[755], c[755]);
HA HA_134(r[661], c[755], r[756], c[756]);
HA HA_135(r[662], c[756], r[757], c[757]);
HA HA_136(r[663], c[757], r[758], c[758]);
HA HA_137(r[664], c[758], r[759], c[759]);
HA HA_138(r[665], c[759], r[760], c[760]);
HA HA_139(r[564], r[666], r[761], c[761]);
FA FA_622(r[667], r[668], c[761], r[762], c[762]);
FA FA_623(r[566], c[667], c[668], r[763], c[763]);
HA HA_140(r[669], c[762], r[764], c[764]);
FA FA_624(r[567], r[568], c[669], r[765], c[765]);
FA FA_625(c[568], r[569], c[670], r[766], c[766]);
HA HA_141(r[671], c[765], r[767], c[767]);
FA FA_626(c[569], r[570], c[671], r[768], c[768]);
FA FA_627(r[571], r[572], c[672], r[769], c[769]);
FA FA_628(c[572], r[573], c[674], r[770], c[770]);
FA FA_629(c[458], r[459], c[573], r[771], c[771]);
HA HA_142(r[574], c[675], r[772], c[772]);
FA FA_630(c[459], r[460], r[461], r[773], c[773]);
FA FA_631(c[461], r[462], r[463], r[774], c[774]);
HA HA_143(c[575], r[576], r[775], c[775]);
FA FA_632(r[464], r[465], r[466], r[776], c[776]);
FA FA_633(r[467], r[468], c[577], r[777], c[777]);
HA HA_144(r[578], r[579], r[778], c[778]);
FA FA_634(r[470], c[578], c[579], r[779], c[779]);
FA FA_635(c[580], c[581], c[582], r[780], c[780]);
FA FA_636(c[584], r[585], r[586], r[781], c[781]);
FA FA_637(c[585], c[586], c[587], r[782], c[782]);
FA FA_638(c[589], r[590], r[591], r[783], c[783]);
FA FA_639(c[590], c[591], c[592], r[784], c[784]);
FA FA_640(r[593], r[594], r[595], r[785], c[785]);
FA FA_641(c[595], r[596], r[597], r[786], c[786]);
HA HA_145(r[598], c[692], r[787], c[787]);
FA FA_642(r[486], c[596], c[597], r[788], c[788]);
FA FA_643(c[598], r[599], r[600], r[789], c[789]);
HA HA_146(c[694], c[695], r[790], c[790]);
FA FA_644(r[488], r[489], c[599], r[791], c[791]);
FA FA_645(c[600], r[601], r[602], r[792], c[792]);
FA FA_646(r[491], r[492], c[601], r[793], c[793]);
FA FA_647(c[602], r[603], r[604], r[794], c[794]);
HA HA_147(c[700], c[701], r[795], c[795]);
FA FA_648(r[494], r[495], c[603], r[796], c[796]);
FA FA_649(c[604], r[605], r[606], r[797], c[797]);
FA FA_650(c[495], r[496], r[497], r[798], c[798]);
FA FA_651(r[498], c[605], c[606], r[799], c[799]);
FA FA_652(r[500], r[501], c[607], r[800], c[800]);
FA FA_653(c[608], c[609], r[610], r[801], c[801]);
HA HA_148(r[611], c[709], r[802], c[802]);
FA FA_654(c[501], r[502], r[503], r[803], c[803]);
FA FA_655(r[504], c[610], c[611], r[804], c[804]);
HA HA_149(r[612], r[613], r[805], c[805]);
FA FA_656(r[506], r[507], c[612], r[806], c[806]);
FA FA_657(c[613], c[614], r[615], r[807], c[807]);
FA FA_658(r[510], c[615], c[616], r[808], c[808]);
FA FA_659(r[617], r[618], r[619], r[809], c[809]);
FA FA_660(c[510], r[511], r[512], r[810], c[810]);
FA FA_661(c[617], c[618], c[619], r[811], c[811]);
HA HA_150(r[620], r[621], r[812], c[812]);
FA FA_662(c[621], r[622], r[623], r[813], c[813]);
FA FA_663(r[624], c[721], c[722], r[814], c[814]);
FA FA_664(r[517], c[622], c[623], r[815], c[815]);
FA FA_665(c[624], r[625], r[626], r[816], c[816]);
HA HA_151(c[723], c[724], r[817], c[817]);
FA FA_666(r[518], r[519], c[625], r[818], c[818]);
FA FA_667(c[626], r[627], r[628], r[819], c[819]);
HA HA_152(c[726], c[727], r[820], c[820]);
FA FA_668(c[628], r[629], r[630], r[821], c[821]);
HA HA_153(r[631], c[729], r[822], c[822]);
FA FA_669(c[629], c[630], c[631], r[823], c[823]);
HA HA_154(r[632], r[633], r[824], c[824]);
FA FA_670(c[633], r[634], r[635], r[825], c[825]);
FA FA_671(c[636], r[637], r[638], r[826], c[826]);
FA FA_672(c[637], c[638], c[639], r[827], c[827]);
FA FA_673(r[534], r[535], c[640], r[828], c[828]);
FA FA_674(r[537], c[642], c[643], r[829], c[829]);
HA HA_155(r[644], r[645], r[830], c[830]);
FA FA_675(r[540], c[644], c[645], r[831], c[831]);
FA FA_676(r[541], r[542], c[646], r[832], c[832]);
HA HA_156(c[647], r[648], r[833], c[833]);
FA FA_677(c[648], r[649], c[743], r[834], c[834]);
FA FA_678(c[544], r[545], c[649], r[835], c[835]);
HA HA_157(r[650], c[744], r[836], c[836]);
FA FA_679(r[651], r[652], c[746], r[837], c[837]);
FA FA_680(c[652], r[653], c[747], r[838], c[838]);
HA HA_158(r[748], c[837], r[839], c[839]);
FA FA_681(r[654], r[655], c[748], r[840], c[840]);
FA FA_682(c[655], r[656], c[749], r[841], c[841]);
HA HA_159(r[750], c[840], r[842], c[842]);
FA FA_683(r[751], r[752], c[841], r[843], c[843]);
HA HA_160(r[753], c[843], r[844], c[844]);
HA HA_161(r[754], c[844], r[845], c[845]);
HA HA_162(r[755], c[845], r[846], c[846]);
HA HA_163(r[756], c[846], r[847], c[847]);
HA HA_164(r[757], c[847], r[848], c[848]);
HA HA_165(r[758], c[848], r[849], c[849]);
HA HA_166(r[759], c[849], r[850], c[850]);
HA HA_167(r[760], c[850], r[851], c[851]);
HA HA_168(r[763], r[764], r[852], c[852]);
FA FA_684(r[670], c[763], c[764], r[853], c[853]);
HA HA_169(r[765], c[852], r[854], c[854]);
FA FA_685(r[766], r[767], c[853], r[855], c[855]);
FA FA_686(r[672], r[673], c[766], r[856], c[856]);
FA FA_687(c[673], r[674], c[768], r[857], c[857]);
HA HA_170(r[769], c[856], r[858], c[858]);
FA FA_688(r[675], r[676], c[769], r[859], c[859]);
FA FA_689(c[676], r[677], c[770], r[860], c[860]);
FA FA_690(c[574], r[575], c[677], r[861], c[861]);
HA HA_171(r[678], c[771], r[862], c[862]);
FA FA_691(c[678], r[679], c[773], r[863], c[863]);
FA FA_692(c[576], r[577], c[679], r[864], c[864]);
HA HA_172(r[680], c[774], r[865], c[865]);
FA FA_693(c[680], r[681], c[776], r[866], c[866]);
FA FA_694(r[580], r[581], r[582], r[867], c[867]);
FA FA_695(r[583], r[584], c[682], r[868], c[868]);
HA HA_173(r[683], r[684], r[869], c[869]);
FA FA_696(r[587], c[683], c[684], r[870], c[870]);
FA FA_697(r[588], r[589], c[685], r[871], c[871]);
FA FA_698(r[592], c[687], c[688], r[872], c[872]);
FA FA_699(c[689], c[690], c[691], r[873], c[873]);
FA FA_700(c[693], r[694], r[695], r[874], c[874]);
FA FA_701(c[696], r[697], r[698], r[875], c[875]);
FA FA_702(c[697], c[698], c[699], r[876], c[876]);
FA FA_703(r[700], r[701], r[702], r[877], c[877]);
FA FA_704(c[702], r[703], r[704], r[878], c[878]);
HA HA_174(r[705], c[791], r[879], c[879]);
FA FA_705(c[703], c[704], c[705], r[880], c[880]);
FA FA_706(r[706], r[707], r[708], r[881], c[881]);
FA FA_707(r[607], r[608], r[609], r[882], c[882]);
FA FA_708(c[706], c[707], c[708], r[883], c[883]);
HA HA_175(r[709], r[710], r[884], c[884]);
FA FA_709(c[710], r[711], r[712], r[885], c[885]);
FA FA_710(r[713], c[798], c[799], r[886], c[886]);
FA FA_711(r[614], c[711], c[712], r[887], c[887]);
FA FA_712(c[713], r[714], r[715], r[888], c[888]);
HA HA_176(c[800], c[801], r[889], c[889]);
FA FA_713(r[616], c[714], c[715], r[890], c[890]);
FA FA_714(r[716], r[717], r[718], r[891], c[891]);
HA HA_177(c[803], c[804], r[892], c[892]);
FA FA_715(c[716], c[717], c[718], r[893], c[893]);
FA FA_716(r[719], r[720], c[806], r[894], c[894]);
FA FA_717(c[719], c[720], r[721], r[895], c[895]);
HA HA_178(r[722], c[808], r[896], c[896]);
FA FA_718(r[723], r[724], r[725], r[897], c[897]);
FA FA_719(c[725], r[726], r[727], r[898], c[898]);
FA FA_720(c[728], r[729], r[730], r[899], c[899]);
FA FA_721(c[730], r[731], r[732], r[900], c[900]);
FA FA_722(c[731], c[732], r[733], r[901], c[901]);
FA FA_723(r[636], c[733], c[734], r[902], c[902]);
FA FA_724(r[639], c[735], c[736], r[903], c[903]);
HA HA_179(r[737], r[738], r[904], c[904]);
FA FA_725(r[640], r[641], c[737], r[905], c[905]);
FA FA_726(c[641], r[642], r[643], r[906], c[906]);
HA HA_180(c[739], r[740], r[907], c[907]);
FA FA_727(c[740], r[741], c[828], r[908], c[908]);
FA FA_728(r[646], r[647], c[741], r[909], c[909]);
HA HA_181(r[742], c[829], r[910], c[910]);
FA FA_729(c[742], r[743], c[831], r[911], c[911]);
FA FA_730(r[744], r[745], c[832], r[912], c[912]);
FA FA_731(c[745], r[746], c[834], r[913], c[913]);
FA FA_732(r[747], c[835], c[836], r[914], c[914]);
HA HA_182(r[837], c[913], r[915], c[915]);
FA FA_733(r[838], r[839], c[914], r[916], c[916]);
FA FA_734(r[749], c[838], c[839], r[917], c[917]);
HA HA_183(r[840], c[916], r[918], c[918]);
FA FA_735(r[841], r[842], c[917], r[919], c[919]);
FA FA_736(c[842], r[843], c[919], r[920], c[920]);
HA HA_184(r[844], c[920], r[921], c[921]);
HA HA_185(r[845], c[921], r[922], c[922]);
HA HA_186(r[846], c[922], r[923], c[923]);
HA HA_187(r[847], c[923], r[924], c[924]);
HA HA_188(r[848], c[924], r[925], c[925]);
HA HA_189(r[849], c[925], r[926], c[926]);
HA HA_190(r[850], c[926], r[927], c[927]);
HA HA_191(r[851], c[927], r[928], c[928]);
HA HA_192(r[853], r[854], r[929], c[929]);
FA FA_737(c[854], r[855], c[929], r[930], c[930]);
FA FA_738(c[767], r[768], c[855], r[931], c[931]);
HA HA_193(r[856], c[930], r[932], c[932]);
FA FA_739(r[857], r[858], c[931], r[933], c[933]);
FA FA_740(r[770], c[857], c[858], r[934], c[934]);
HA HA_194(r[859], c[933], r[935], c[935]);
FA FA_741(r[771], r[772], c[859], r[936], c[936]);
FA FA_742(c[772], r[773], c[860], r[937], c[937]);
FA FA_743(r[774], r[775], c[861], r[938], c[938]);
FA FA_744(c[775], r[776], c[863], r[939], c[939]);
FA FA_745(r[777], r[778], c[864], r[940], c[940]);
FA FA_746(c[681], r[682], c[777], r[941], c[941]);
HA HA_195(c[778], r[779], r[942], c[942]);
FA FA_747(c[779], r[780], c[867], r[943], c[943]);
FA FA_748(r[685], r[686], c[780], r[944], c[944]);
HA HA_196(r[781], c[868], r[945], c[945]);
FA FA_749(c[686], r[687], r[688], r[946], c[946]);
FA FA_750(r[689], r[690], r[691], r[947], c[947]);
HA HA_197(c[782], r[783], r[948], c[948]);
FA FA_751(r[692], r[693], c[783], r[949], c[949]);
FA FA_752(r[696], c[784], c[785], r[950], c[950]);
HA HA_198(r[786], r[787], r[951], c[951]);
FA FA_753(r[699], c[786], c[787], r[952], c[952]);
FA FA_754(c[788], c[789], c[790], r[953], c[953]);
FA FA_755(c[792], r[793], r[794], r[954], c[954]);
FA FA_756(c[793], c[794], c[795], r[955], c[955]);
FA FA_757(c[796], c[797], r[798], r[956], c[956]);
FA FA_758(r[800], r[801], r[802], r[957], c[957]);
FA FA_759(c[802], r[803], r[804], r[958], c[958]);
FA FA_760(c[805], r[806], r[807], r[959], c[959]);
FA FA_761(c[807], r[808], r[809], r[960], c[960]);
FA FA_762(c[809], r[810], r[811], r[961], c[961]);
FA FA_763(c[810], c[811], c[812], r[962], c[962]);
FA FA_764(r[728], c[813], c[814], r[963], c[963]);
FA FA_765(c[815], c[816], c[817], r[964], c[964]);
FA FA_766(c[818], c[819], c[820], r[965], c[965]);
HA HA_199(r[821], r[822], r[966], c[966]);
FA FA_767(r[734], c[821], c[822], r[967], c[967]);
FA FA_768(r[735], r[736], c[823], r[968], c[968]);
HA HA_200(c[824], r[825], r[969], c[969]);
FA FA_769(c[825], r[826], c[902], r[970], c[970]);
FA FA_770(c[738], r[739], c[826], r[971], c[971]);
HA HA_201(r[827], c[903], r[972], c[972]);
FA FA_771(c[827], r[828], c[905], r[973], c[973]);
FA FA_772(r[829], r[830], c[906], r[974], c[974]);
FA FA_773(c[830], r[831], c[908], r[975], c[975]);
FA FA_774(r[832], r[833], c[909], r[976], c[976]);
FA FA_775(c[833], r[834], c[911], r[977], c[977]);
HA HA_202(r[912], c[976], r[978], c[978]);
FA FA_776(r[835], r[836], c[912], r[979], c[979]);
FA FA_777(r[914], r[915], c[979], r[980], c[980]);
FA FA_778(c[915], r[916], c[980], r[981], c[981]);
FA FA_779(r[917], r[918], c[981], r[982], c[982]);
FA FA_780(c[918], r[919], c[982], r[983], c[983]);
HA HA_203(r[920], c[983], r[984], c[984]);
HA HA_204(r[921], c[984], r[985], c[985]);
HA HA_205(r[922], c[985], r[986], c[986]);
HA HA_206(r[923], c[986], r[987], c[987]);
HA HA_207(r[924], c[987], r[988], c[988]);
HA HA_208(r[925], c[988], r[989], c[989]);
HA HA_209(r[926], c[989], r[990], c[990]);
HA HA_210(r[927], c[990], r[991], c[991]);
HA HA_211(r[928], c[991], r[992], c[992]);
HA HA_212(r[931], r[932], r[993], c[993]);
FA FA_781(c[932], r[933], c[993], r[994], c[994]);
FA FA_782(r[934], r[935], c[994], r[995], c[995]);
FA FA_783(r[860], c[934], c[935], r[996], c[996]);
HA HA_213(r[936], c[995], r[997], c[997]);
FA FA_784(r[861], r[862], c[936], r[998], c[998]);
FA FA_785(c[862], r[863], c[937], r[999], c[999]);
HA HA_214(r[938], c[998], r[1000], c[1000]);
FA FA_786(r[864], r[865], c[938], r[1001], c[1001]);
FA FA_787(c[865], r[866], c[939], r[1002], c[1002]);
HA HA_215(r[940], c[1001], r[1003], c[1003]);
FA FA_788(c[866], r[867], c[940], r[1004], c[1004]);
FA FA_789(r[868], r[869], c[941], r[1005], c[1005]);
FA FA_790(c[869], r[870], c[943], r[1006], c[1006]);
FA FA_791(c[781], r[782], c[870], r[1007], c[1007]);
HA HA_216(r[871], c[944], r[1008], c[1008]);
FA FA_792(c[871], r[872], c[946], r[1009], c[1009]);
FA FA_793(r[784], r[785], c[872], r[1010], c[1010]);
HA HA_217(r[873], c[947], r[1011], c[1011]);
FA FA_794(c[873], r[874], c[949], r[1012], c[1012]);
FA FA_795(r[788], r[789], r[790], r[1013], c[1013]);
FA FA_796(r[791], r[792], c[875], r[1014], c[1014]);
HA HA_218(r[876], r[877], r[1015], c[1015]);
FA FA_797(r[795], c[876], c[877], r[1016], c[1016]);
FA FA_798(r[796], r[797], c[878], r[1017], c[1017]);
FA FA_799(r[799], c[880], c[881], r[1018], c[1018]);
FA FA_800(c[882], c[883], c[884], r[1019], c[1019]);
HA HA_219(r[885], r[886], r[1020], c[1020]);
FA FA_801(r[805], c[885], c[886], r[1021], c[1021]);
FA FA_802(c[887], c[888], c[889], r[1022], c[1022]);
FA FA_803(c[890], c[891], c[892], r[1023], c[1023]);
HA HA_220(r[893], r[894], r[1024], c[1024]);
FA FA_804(r[812], c[893], c[894], r[1025], c[1025]);
FA FA_805(r[813], r[814], c[895], r[1026], c[1026]);
HA HA_221(c[896], r[897], r[1027], c[1027]);
FA FA_806(r[815], r[816], r[817], r[1028], c[1028]);
FA FA_807(r[818], r[819], r[820], r[1029], c[1029]);
HA HA_222(c[898], r[899], r[1030], c[1030]);
FA FA_808(c[899], r[900], c[964], r[1031], c[1031]);
FA FA_809(r[823], r[824], c[900], r[1032], c[1032]);
HA HA_223(r[901], c[965], r[1033], c[1033]);
FA FA_810(c[901], r[902], c[967], r[1034], c[1034]);
FA FA_811(r[903], r[904], c[968], r[1035], c[1035]);
FA FA_812(c[904], r[905], c[970], r[1036], c[1036]);
FA FA_813(r[906], r[907], c[971], r[1037], c[1037]);
FA FA_814(c[907], r[908], c[973], r[1038], c[1038]);
HA HA_224(r[974], c[1037], r[1039], c[1039]);
FA FA_815(r[909], r[910], c[974], r[1040], c[1040]);
FA FA_816(c[910], r[911], c[975], r[1041], c[1041]);
HA HA_225(r[976], c[1040], r[1042], c[1042]);
FA FA_817(r[977], r[978], c[1041], r[1043], c[1043]);
FA FA_818(r[913], c[977], c[978], r[1044], c[1044]);
HA HA_226(r[979], c[1043], r[1045], c[1045]);
FA FA_819(r[980], c[1044], c[1045], r[1046], c[1046]);
HA HA_227(r[981], c[1046], r[1047], c[1047]);
HA HA_228(r[982], c[1047], r[1048], c[1048]);
HA HA_229(r[983], c[1048], r[1049], c[1049]);
HA HA_230(r[984], c[1049], r[1050], c[1050]);
HA HA_231(r[985], c[1050], r[1051], c[1051]);
HA HA_232(r[986], c[1051], r[1052], c[1052]);
HA HA_233(r[987], c[1052], r[1053], c[1053]);
HA HA_234(r[988], c[1053], r[1054], c[1054]);
HA HA_235(r[989], c[1054], r[1055], c[1055]);
HA HA_236(r[990], c[1055], r[1056], c[1056]);
HA HA_237(r[991], c[1056], r[1057], c[1057]);
HA HA_238(r[992], c[1057], r[1058], c[1058]);
HA HA_239(r[996], r[997], r[1059], c[1059]);
FA FA_820(r[937], c[996], c[997], r[1060], c[1060]);
HA HA_240(r[998], c[1059], r[1061], c[1061]);
FA FA_821(r[999], r[1000], c[1060], r[1062], c[1062]);
FA FA_822(r[939], c[999], c[1000], r[1063], c[1063]);
HA HA_241(r[1001], c[1062], r[1064], c[1064]);
FA FA_823(r[1002], r[1003], c[1063], r[1065], c[1065]);
FA FA_824(r[941], r[942], c[1002], r[1066], c[1066]);
FA FA_825(c[942], r[943], c[1004], r[1067], c[1067]);
HA HA_242(r[1005], c[1066], r[1068], c[1068]);
FA FA_826(r[944], r[945], c[1005], r[1069], c[1069]);
FA FA_827(c[945], r[946], c[1006], r[1070], c[1070]);
FA FA_828(r[947], r[948], c[1007], r[1071], c[1071]);
FA FA_829(c[948], r[949], c[1009], r[1072], c[1072]);
FA FA_830(r[950], r[951], c[1010], r[1073], c[1073]);
FA FA_831(c[874], r[875], c[950], r[1074], c[1074]);
HA HA_243(c[951], r[952], r[1075], c[1075]);
FA FA_832(c[952], r[953], c[1013], r[1076], c[1076]);
FA FA_833(r[878], r[879], c[953], r[1077], c[1077]);
HA HA_244(r[954], c[1014], r[1078], c[1078]);
FA FA_834(c[879], r[880], r[881], r[1079], c[1079]);
FA FA_835(r[882], r[883], r[884], r[1080], c[1080]);
HA HA_245(c[955], r[956], r[1081], c[1081]);
FA FA_836(c[956], r[957], c[1018], r[1082], c[1082]);
FA FA_837(r[887], r[888], r[889], r[1083], c[1083]);
FA FA_838(r[890], r[891], r[892], r[1084], c[1084]);
HA HA_246(c[958], r[959], r[1085], c[1085]);
FA FA_839(c[959], r[960], c[1022], r[1086], c[1086]);
FA FA_840(r[895], r[896], c[960], r[1087], c[1087]);
HA HA_247(r[961], c[1023], r[1088], c[1088]);
FA FA_841(c[961], r[962], c[1025], r[1089], c[1089]);
FA FA_842(c[897], r[898], c[962], r[1090], c[1090]);
HA HA_248(r[963], c[1026], r[1091], c[1091]);
FA FA_843(c[963], r[964], c[1028], r[1092], c[1092]);
FA FA_844(r[965], r[966], c[1029], r[1093], c[1093]);
FA FA_845(c[966], r[967], c[1031], r[1094], c[1094]);
FA FA_846(r[968], r[969], c[1032], r[1095], c[1095]);
FA FA_847(c[969], r[970], c[1034], r[1096], c[1096]);
HA HA_249(r[1035], c[1095], r[1097], c[1097]);
FA FA_848(r[971], r[972], c[1035], r[1098], c[1098]);
FA FA_849(c[972], r[973], c[1036], r[1099], c[1099]);
HA HA_250(r[1037], c[1098], r[1100], c[1100]);
FA FA_850(r[1038], r[1039], c[1099], r[1101], c[1101]);
FA FA_851(r[975], c[1038], c[1039], r[1102], c[1102]);
HA HA_251(r[1040], c[1101], r[1103], c[1103]);
FA FA_852(r[1041], r[1042], c[1102], r[1104], c[1104]);
FA FA_853(c[1042], r[1043], c[1104], r[1105], c[1105]);
FA FA_854(r[1044], r[1045], c[1105], r[1106], c[1106]);
HA HA_252(r[1046], c[1106], r[1107], c[1107]);
HA HA_253(r[1047], c[1107], r[1108], c[1108]);
HA HA_254(r[1048], c[1108], r[1109], c[1109]);
HA HA_255(r[1049], c[1109], r[1110], c[1110]);
HA HA_256(r[1050], c[1110], r[1111], c[1111]);
HA HA_257(r[1051], c[1111], r[1112], c[1112]);
HA HA_258(r[1052], c[1112], r[1113], c[1113]);
HA HA_259(r[1053], c[1113], r[1114], c[1114]);
HA HA_260(r[1054], c[1114], r[1115], c[1115]);
HA HA_261(r[1055], c[1115], r[1116], c[1116]);
HA HA_262(r[1056], c[1116], r[1117], c[1117]);
HA HA_263(r[1057], c[1117], r[1118], c[1118]);
HA HA_264(r[1058], c[1118], r[1119], c[1119]);
HA HA_265(r[1060], r[1061], r[1120], c[1120]);
FA FA_855(c[1061], r[1062], c[1120], r[1121], c[1121]);
FA FA_856(r[1063], r[1064], c[1121], r[1122], c[1122]);
FA FA_857(c[1064], r[1065], c[1122], r[1123], c[1123]);
FA FA_858(c[1003], r[1004], c[1065], r[1124], c[1124]);
HA HA_266(r[1066], c[1123], r[1125], c[1125]);
FA FA_859(r[1067], r[1068], c[1124], r[1126], c[1126]);
FA FA_860(r[1006], c[1067], c[1068], r[1127], c[1127]);
HA HA_267(r[1069], c[1126], r[1128], c[1128]);
FA FA_861(r[1007], r[1008], c[1069], r[1129], c[1129]);
FA FA_862(c[1008], r[1009], c[1070], r[1130], c[1130]);
HA HA_268(r[1071], c[1129], r[1131], c[1131]);
FA FA_863(r[1010], r[1011], c[1071], r[1132], c[1132]);
FA FA_864(c[1011], r[1012], c[1072], r[1133], c[1133]);
HA HA_269(r[1073], c[1132], r[1134], c[1134]);
FA FA_865(c[1012], r[1013], c[1073], r[1135], c[1135]);
FA FA_866(r[1014], r[1015], c[1074], r[1136], c[1136]);
FA FA_867(c[1015], r[1016], c[1076], r[1137], c[1137]);
FA FA_868(c[954], r[955], c[1016], r[1138], c[1138]);
HA HA_270(r[1017], c[1077], r[1139], c[1139]);
FA FA_869(c[1017], r[1018], c[1079], r[1140], c[1140]);
FA FA_870(r[1019], r[1020], c[1080], r[1141], c[1141]);
FA FA_871(c[957], r[958], c[1019], r[1142], c[1142]);
HA HA_271(c[1020], r[1021], r[1143], c[1143]);
FA FA_872(c[1021], r[1022], c[1083], r[1144], c[1144]);
FA FA_873(r[1023], r[1024], c[1084], r[1145], c[1145]);
FA FA_874(c[1024], r[1025], c[1086], r[1146], c[1146]);
FA FA_875(r[1026], r[1027], c[1087], r[1147], c[1147]);
FA FA_876(c[1027], r[1028], c[1089], r[1148], c[1148]);
FA FA_877(r[1029], r[1030], c[1090], r[1149], c[1149]);
FA FA_878(c[1030], r[1031], c[1092], r[1150], c[1150]);
HA HA_272(r[1093], c[1149], r[1151], c[1151]);
FA FA_879(r[1032], r[1033], c[1093], r[1152], c[1152]);
FA FA_880(c[1033], r[1034], c[1094], r[1153], c[1153]);
HA HA_273(r[1095], c[1152], r[1154], c[1154]);
FA FA_881(r[1096], r[1097], c[1153], r[1155], c[1155]);
FA FA_882(r[1036], c[1096], c[1097], r[1156], c[1156]);
HA HA_274(r[1098], c[1155], r[1157], c[1157]);
FA FA_883(r[1099], r[1100], c[1156], r[1158], c[1158]);
FA FA_884(c[1100], r[1101], c[1158], r[1159], c[1159]);
FA FA_885(r[1102], r[1103], c[1159], r[1160], c[1160]);
FA FA_886(c[1103], r[1104], c[1160], r[1161], c[1161]);
HA HA_275(r[1105], c[1161], r[1162], c[1162]);
HA HA_276(r[1106], c[1162], r[1163], c[1163]);
HA HA_277(r[1107], c[1163], r[1164], c[1164]);
HA HA_278(r[1108], c[1164], r[1165], c[1165]);
HA HA_279(r[1109], c[1165], r[1166], c[1166]);
HA HA_280(r[1110], c[1166], r[1167], c[1167]);
HA HA_281(r[1111], c[1167], r[1168], c[1168]);
HA HA_282(r[1112], c[1168], r[1169], c[1169]);
HA HA_283(r[1113], c[1169], r[1170], c[1170]);
HA HA_284(r[1114], c[1170], r[1171], c[1171]);
HA HA_285(r[1115], c[1171], r[1172], c[1172]);
HA HA_286(r[1116], c[1172], r[1173], c[1173]);
HA HA_287(r[1117], c[1173], r[1174], c[1174]);
HA HA_288(r[1118], c[1174], r[1175], c[1175]);
HA HA_289(r[1119], c[1175], r[1176], c[1176]);
HA HA_290(r[1124], r[1125], r[1177], c[1177]);
FA FA_887(c[1125], r[1126], c[1177], r[1178], c[1178]);
FA FA_888(r[1127], r[1128], c[1178], r[1179], c[1179]);
FA FA_889(r[1070], c[1127], c[1128], r[1180], c[1180]);
HA HA_291(r[1129], c[1179], r[1181], c[1181]);
FA FA_890(r[1130], r[1131], c[1180], r[1182], c[1182]);
FA FA_891(r[1072], c[1130], c[1131], r[1183], c[1183]);
HA HA_292(r[1132], c[1182], r[1184], c[1184]);
FA FA_892(r[1133], r[1134], c[1183], r[1185], c[1185]);
FA FA_893(r[1074], r[1075], c[1133], r[1186], c[1186]);
FA FA_894(c[1075], r[1076], c[1135], r[1187], c[1187]);
HA HA_293(r[1136], c[1186], r[1188], c[1188]);
FA FA_895(r[1077], r[1078], c[1136], r[1189], c[1189]);
FA FA_896(c[1078], r[1079], c[1137], r[1190], c[1190]);
FA FA_897(r[1080], r[1081], c[1138], r[1191], c[1191]);
FA FA_898(c[1081], r[1082], c[1140], r[1192], c[1192]);
HA HA_294(r[1141], c[1191], r[1193], c[1193]);
FA FA_899(c[1082], r[1083], c[1141], r[1194], c[1194]);
FA FA_900(r[1084], r[1085], c[1142], r[1195], c[1195]);
FA FA_901(c[1085], r[1086], c[1144], r[1196], c[1196]);
HA HA_295(r[1145], c[1195], r[1197], c[1197]);
FA FA_902(r[1087], r[1088], c[1145], r[1198], c[1198]);
FA FA_903(c[1088], r[1089], c[1146], r[1199], c[1199]);
HA HA_296(r[1147], c[1198], r[1200], c[1200]);
FA FA_904(r[1090], r[1091], c[1147], r[1201], c[1201]);
FA FA_905(c[1091], r[1092], c[1148], r[1202], c[1202]);
HA HA_297(r[1149], c[1201], r[1203], c[1203]);
FA FA_906(r[1150], r[1151], c[1202], r[1204], c[1204]);
FA FA_907(r[1094], c[1150], c[1151], r[1205], c[1205]);
HA HA_298(r[1152], c[1204], r[1206], c[1206]);
FA FA_908(r[1153], r[1154], c[1205], r[1207], c[1207]);
FA FA_909(c[1154], r[1155], c[1207], r[1208], c[1208]);
FA FA_910(r[1156], r[1157], c[1208], r[1209], c[1209]);
FA FA_911(c[1157], r[1158], c[1209], r[1210], c[1210]);
HA HA_299(r[1159], c[1210], r[1211], c[1211]);
HA HA_300(r[1160], c[1211], r[1212], c[1212]);
HA HA_301(r[1161], c[1212], r[1213], c[1213]);
HA HA_302(r[1162], c[1213], r[1214], c[1214]);
HA HA_303(r[1163], c[1214], r[1215], c[1215]);
HA HA_304(r[1164], c[1215], r[1216], c[1216]);
HA HA_305(r[1165], c[1216], r[1217], c[1217]);
HA HA_306(r[1166], c[1217], r[1218], c[1218]);
HA HA_307(r[1167], c[1218], r[1219], c[1219]);
HA HA_308(r[1168], c[1219], r[1220], c[1220]);
HA HA_309(r[1169], c[1220], r[1221], c[1221]);
HA HA_310(r[1170], c[1221], r[1222], c[1222]);
HA HA_311(r[1171], c[1222], r[1223], c[1223]);
HA HA_312(r[1172], c[1223], r[1224], c[1224]);
HA HA_313(r[1173], c[1224], r[1225], c[1225]);
HA HA_314(r[1174], c[1225], r[1226], c[1226]);
HA HA_315(r[1175], c[1226], r[1227], c[1227]);
HA HA_316(r[1176], c[1227], r[1228], c[1228]);
HA HA_317(r[1180], r[1181], r[1229], c[1229]);
FA FA_912(c[1181], r[1182], c[1229], r[1230], c[1230]);
FA FA_913(r[1183], r[1184], c[1230], r[1231], c[1231]);
FA FA_914(c[1184], r[1185], c[1231], r[1232], c[1232]);
FA FA_915(c[1134], r[1135], c[1185], r[1233], c[1233]);
HA HA_318(r[1186], c[1232], r[1234], c[1234]);
FA FA_916(r[1187], r[1188], c[1233], r[1235], c[1235]);
FA FA_917(r[1137], c[1187], c[1188], r[1236], c[1236]);
HA HA_319(r[1189], c[1235], r[1237], c[1237]);
FA FA_918(r[1138], r[1139], c[1189], r[1238], c[1238]);
FA FA_919(c[1139], r[1140], c[1190], r[1239], c[1239]);
HA HA_320(r[1191], c[1238], r[1240], c[1240]);
FA FA_920(r[1192], r[1193], c[1239], r[1241], c[1241]);
FA FA_921(r[1142], r[1143], c[1192], r[1242], c[1242]);
FA FA_922(c[1143], r[1144], c[1194], r[1243], c[1243]);
HA HA_321(r[1195], c[1242], r[1244], c[1244]);
FA FA_923(r[1196], r[1197], c[1243], r[1245], c[1245]);
FA FA_924(r[1146], c[1196], c[1197], r[1246], c[1246]);
HA HA_322(r[1198], c[1245], r[1247], c[1247]);
FA FA_925(r[1199], r[1200], c[1246], r[1248], c[1248]);
FA FA_926(r[1148], c[1199], c[1200], r[1249], c[1249]);
HA HA_323(r[1201], c[1248], r[1250], c[1250]);
FA FA_927(r[1202], r[1203], c[1249], r[1251], c[1251]);
FA FA_928(c[1203], r[1204], c[1251], r[1252], c[1252]);
FA FA_929(r[1205], r[1206], c[1252], r[1253], c[1253]);
FA FA_930(c[1206], r[1207], c[1253], r[1254], c[1254]);
HA HA_324(r[1208], c[1254], r[1255], c[1255]);
HA HA_325(r[1209], c[1255], r[1256], c[1256]);
HA HA_326(r[1210], c[1256], r[1257], c[1257]);
HA HA_327(r[1211], c[1257], r[1258], c[1258]);
HA HA_328(r[1212], c[1258], r[1259], c[1259]);
HA HA_329(r[1213], c[1259], r[1260], c[1260]);
HA HA_330(r[1214], c[1260], r[1261], c[1261]);
HA HA_331(r[1215], c[1261], r[1262], c[1262]);
HA HA_332(r[1216], c[1262], r[1263], c[1263]);
HA HA_333(r[1217], c[1263], r[1264], c[1264]);
HA HA_334(r[1218], c[1264], r[1265], c[1265]);
HA HA_335(r[1219], c[1265], r[1266], c[1266]);
HA HA_336(r[1220], c[1266], r[1267], c[1267]);
HA HA_337(r[1221], c[1267], r[1268], c[1268]);
HA HA_338(r[1222], c[1268], r[1269], c[1269]);
HA HA_339(r[1223], c[1269], r[1270], c[1270]);
HA HA_340(r[1224], c[1270], r[1271], c[1271]);
HA HA_341(r[1225], c[1271], r[1272], c[1272]);
HA HA_342(r[1226], c[1272], r[1273], c[1273]);
HA HA_343(r[1227], c[1273], r[1274], c[1274]);
HA HA_344(r[1228], c[1274], r[1275], c[1275]);
HA HA_345(r[1233], r[1234], r[1276], c[1276]);
FA FA_931(c[1234], r[1235], c[1276], r[1277], c[1277]);
FA FA_932(r[1236], r[1237], c[1277], r[1278], c[1278]);
FA FA_933(r[1190], c[1236], c[1237], r[1279], c[1279]);
HA HA_346(r[1238], c[1278], r[1280], c[1280]);
FA FA_934(r[1239], r[1240], c[1279], r[1281], c[1281]);
FA FA_935(c[1240], r[1241], c[1281], r[1282], c[1282]);
FA FA_936(c[1193], r[1194], c[1241], r[1283], c[1283]);
HA HA_347(r[1242], c[1282], r[1284], c[1284]);
FA FA_937(r[1243], r[1244], c[1283], r[1285], c[1285]);
FA FA_938(c[1244], r[1245], c[1285], r[1286], c[1286]);
FA FA_939(r[1246], r[1247], c[1286], r[1287], c[1287]);
FA FA_940(c[1247], r[1248], c[1287], r[1288], c[1288]);
FA FA_941(r[1249], r[1250], c[1288], r[1289], c[1289]);
FA FA_942(c[1250], r[1251], c[1289], r[1290], c[1290]);
HA HA_348(r[1252], c[1290], r[1291], c[1291]);
HA HA_349(r[1253], c[1291], r[1292], c[1292]);
HA HA_350(r[1254], c[1292], r[1293], c[1293]);
HA HA_351(r[1255], c[1293], r[1294], c[1294]);
HA HA_352(r[1256], c[1294], r[1295], c[1295]);
HA HA_353(r[1257], c[1295], r[1296], c[1296]);
HA HA_354(r[1258], c[1296], r[1297], c[1297]);
HA HA_355(r[1259], c[1297], r[1298], c[1298]);
HA HA_356(r[1260], c[1298], r[1299], c[1299]);
HA HA_357(r[1261], c[1299], r[1300], c[1300]);
HA HA_358(r[1262], c[1300], r[1301], c[1301]);
HA HA_359(r[1263], c[1301], r[1302], c[1302]);
HA HA_360(r[1264], c[1302], r[1303], c[1303]);
HA HA_361(r[1265], c[1303], r[1304], c[1304]);
HA HA_362(r[1266], c[1304], r[1305], c[1305]);
HA HA_363(r[1267], c[1305], r[1306], c[1306]);
HA HA_364(r[1268], c[1306], r[1307], c[1307]);
HA HA_365(r[1269], c[1307], r[1308], c[1308]);
HA HA_366(r[1270], c[1308], r[1309], c[1309]);
HA HA_367(r[1271], c[1309], r[1310], c[1310]);
HA HA_368(r[1272], c[1310], r[1311], c[1311]);
HA HA_369(r[1273], c[1311], r[1312], c[1312]);
HA HA_370(r[1274], c[1312], r[1313], c[1313]);
HA HA_371(r[1275], c[1313], r[1314], c[1314]);
HA HA_372(r[1279], r[1280], r[1315], c[1315]);
FA FA_943(c[1280], r[1281], c[1315], r[1316], c[1316]);
HA HA_373(r[1282], c[1316], r[1317], c[1317]);
FA FA_944(r[1283], r[1284], c[1317], r[1318], c[1318]);
FA FA_945(c[1284], r[1285], c[1318], r[1319], c[1319]);
HA HA_374(r[1286], c[1319], r[1320], c[1320]);
HA HA_375(r[1287], c[1320], r[1321], c[1321]);
HA HA_376(r[1288], c[1321], r[1322], c[1322]);
HA HA_377(r[1289], c[1322], r[1323], c[1323]);
HA HA_378(r[1290], c[1323], r[1324], c[1324]);
HA HA_379(r[1291], c[1324], r[1325], c[1325]);
HA HA_380(r[1292], c[1325], r[1326], c[1326]);
HA HA_381(r[1293], c[1326], r[1327], c[1327]);
HA HA_382(r[1294], c[1327], r[1328], c[1328]);
HA HA_383(r[1295], c[1328], r[1329], c[1329]);
HA HA_384(r[1296], c[1329], r[1330], c[1330]);
HA HA_385(r[1297], c[1330], r[1331], c[1331]);
HA HA_386(r[1298], c[1331], r[1332], c[1332]);
HA HA_387(r[1299], c[1332], r[1333], c[1333]);
HA HA_388(r[1300], c[1333], r[1334], c[1334]);
HA HA_389(r[1301], c[1334], r[1335], c[1335]);
HA HA_390(r[1302], c[1335], r[1336], c[1336]);
HA HA_391(r[1303], c[1336], r[1337], c[1337]);
HA HA_392(r[1304], c[1337], r[1338], c[1338]);
HA HA_393(r[1305], c[1338], r[1339], c[1339]);
HA HA_394(r[1306], c[1339], r[1340], c[1340]);
HA HA_395(r[1307], c[1340], r[1341], c[1341]);
HA HA_396(r[1308], c[1341], r[1342], c[1342]);
HA HA_397(r[1309], c[1342], r[1343], c[1343]);
HA HA_398(r[1310], c[1343], r[1344], c[1344]);
HA HA_399(r[1311], c[1344], r[1345], c[1345]);
HA HA_400(r[1312], c[1345], r[1346], c[1346]);
HA HA_401(r[1313], c[1346], r[1347], c[1347]);
HA HA_402(r[1314], c[1347], r[1348], c[1348]);

assign result[0] = p[0][0];
assign result[1] = r[0];
assign result[2] = r[175];
assign result[3] = r[176];
assign result[4] = r[445];
assign result[5] = r[446];
assign result[6] = r[563];
assign result[7] = r[761];
assign result[8] = r[762];
assign result[9] = r[852];
assign result[10] = r[929];
assign result[11] = r[930];
assign result[12] = r[993];
assign result[13] = r[994];
assign result[14] = r[995];
assign result[15] = r[1059];
assign result[16] = r[1120];
assign result[17] = r[1121];
assign result[18] = r[1122];
assign result[19] = r[1123];
assign result[20] = r[1177];
assign result[21] = r[1178];
assign result[22] = r[1179];
assign result[23] = r[1229];
assign result[24] = r[1230];
assign result[25] = r[1231];
assign result[26] = r[1232];
assign result[27] = r[1276];
assign result[28] = r[1277];
assign result[29] = r[1278];
assign result[30] = r[1315];
assign result[31] = r[1316];
assign result[32] = r[1317];
assign result[33] = r[1318];
assign result[34] = r[1319];
assign result[35] = r[1320];
assign result[36] = r[1321];
assign result[37] = r[1322];
assign result[38] = r[1323];
assign result[39] = r[1324];
assign result[40] = r[1325];
assign result[41] = r[1326];
assign result[42] = r[1327];
assign result[43] = r[1328];
assign result[44] = r[1329];
assign result[45] = r[1330];
assign result[46] = r[1331];
assign result[47] = r[1332];
assign result[48] = r[1333];
assign result[49] = r[1334];
assign result[50] = r[1335];
assign result[51] = r[1336];
assign result[52] = r[1337];
assign result[53] = r[1338];
assign result[54] = r[1339];
assign result[55] = r[1340];
assign result[56] = r[1341];
assign result[57] = r[1342];
assign result[58] = r[1343];
assign result[59] = r[1344];
assign result[60] = r[1345];
assign result[61] = r[1346];
assign result[62] = r[1347];
assign result[63] = r[1348];


endmodule

module registerNbits #(
    parameter N = 8
) (
    clk,
    reset,
    en,
    inp,
    out
);
  input clk, reset, en;
  output reg [N-1:0] out;
  input [N-1:0] inp;
  always @(posedge clk) begin
    if (reset) out <= 'b0;
    else if (en) out <= inp;

  end
endmodule


module signed_wallace (
    input i_clk,
    input i_rst,
    input i_en,
    input [31:0] i_inputA,
    input [31:0] i_inputB,
    output [63:0] o_result
);

  wire [31:0] A_reg;
  wire [31:0] B_reg;
  wire [63:0] out_reg;


  registerNbits #(32) regA (
      i_clk,
      i_rst,
      i_en,
      i_inputA,
      A_reg
  );
  registerNbits #(32) regB (
      i_clk,
      i_rst,
      i_en,
      i_inputB,
      B_reg
  );
  signed_wallace_tree_multipler unt (
      A_reg,
      B_reg,
      out_reg
  );
  registerNbits #(64) outReg (
      i_clk,
      i_rst,
      i_en,
      out_reg,
      o_result[63:0]
  );


endmodule