
// 	Tue Dec 20 16:15:44 2022
//	vlsi
//	localhost.localdomain

module registerNbits__parameterized0 (clk_CTS_1_PP_0, clk, reset, en, inp, out);

output [63:0] out;
input clk;
input en;
input [63:0] inp;
input reset;
input clk_CTS_1_PP_0;
wire n_0_0;
wire n_1;
wire CTS_n_tid0_10;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid0_11;
wire hfn_ipo_n6;


AND2_X1 i_0_65 (.ZN (n_65), .A1 (hfn_ipo_n6), .A2 (inp[63]));
AND2_X1 i_0_64 (.ZN (n_64), .A1 (hfn_ipo_n6), .A2 (inp[62]));
AND2_X1 i_0_63 (.ZN (n_63), .A1 (hfn_ipo_n6), .A2 (inp[61]));
AND2_X1 i_0_62 (.ZN (n_62), .A1 (hfn_ipo_n6), .A2 (inp[60]));
AND2_X1 i_0_61 (.ZN (n_61), .A1 (hfn_ipo_n6), .A2 (inp[59]));
AND2_X1 i_0_60 (.ZN (n_60), .A1 (hfn_ipo_n6), .A2 (inp[58]));
AND2_X1 i_0_59 (.ZN (n_59), .A1 (hfn_ipo_n6), .A2 (inp[57]));
AND2_X1 i_0_58 (.ZN (n_58), .A1 (hfn_ipo_n6), .A2 (inp[56]));
AND2_X1 i_0_57 (.ZN (n_57), .A1 (hfn_ipo_n6), .A2 (inp[55]));
AND2_X1 i_0_56 (.ZN (n_56), .A1 (hfn_ipo_n6), .A2 (inp[54]));
AND2_X1 i_0_55 (.ZN (n_55), .A1 (hfn_ipo_n6), .A2 (inp[53]));
AND2_X1 i_0_54 (.ZN (n_54), .A1 (hfn_ipo_n6), .A2 (inp[52]));
AND2_X1 i_0_53 (.ZN (n_53), .A1 (hfn_ipo_n6), .A2 (inp[51]));
AND2_X1 i_0_52 (.ZN (n_52), .A1 (hfn_ipo_n6), .A2 (inp[50]));
AND2_X1 i_0_51 (.ZN (n_51), .A1 (n_0_0), .A2 (inp[49]));
AND2_X1 i_0_50 (.ZN (n_50), .A1 (n_0_0), .A2 (inp[48]));
AND2_X1 i_0_49 (.ZN (n_49), .A1 (n_0_0), .A2 (inp[47]));
AND2_X1 i_0_48 (.ZN (n_48), .A1 (n_0_0), .A2 (inp[46]));
AND2_X1 i_0_47 (.ZN (n_47), .A1 (n_0_0), .A2 (inp[45]));
AND2_X1 i_0_46 (.ZN (n_46), .A1 (n_0_0), .A2 (inp[44]));
AND2_X1 i_0_45 (.ZN (n_45), .A1 (n_0_0), .A2 (inp[43]));
AND2_X1 i_0_44 (.ZN (n_44), .A1 (n_0_0), .A2 (inp[42]));
AND2_X1 i_0_43 (.ZN (n_43), .A1 (n_0_0), .A2 (inp[41]));
AND2_X1 i_0_42 (.ZN (n_42), .A1 (n_0_0), .A2 (inp[40]));
AND2_X1 i_0_41 (.ZN (n_41), .A1 (n_0_0), .A2 (inp[39]));
AND2_X1 i_0_40 (.ZN (n_40), .A1 (n_0_0), .A2 (inp[38]));
AND2_X1 i_0_39 (.ZN (n_39), .A1 (n_0_0), .A2 (inp[37]));
AND2_X1 i_0_38 (.ZN (n_38), .A1 (n_0_0), .A2 (inp[36]));
AND2_X1 i_0_37 (.ZN (n_37), .A1 (n_0_0), .A2 (inp[35]));
AND2_X1 i_0_36 (.ZN (n_36), .A1 (n_0_0), .A2 (inp[34]));
AND2_X1 i_0_35 (.ZN (n_35), .A1 (n_0_0), .A2 (inp[33]));
AND2_X1 i_0_34 (.ZN (n_34), .A1 (n_0_0), .A2 (inp[32]));
AND2_X1 i_0_33 (.ZN (n_33), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (n_32), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (n_31), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (n_30), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (n_29), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (n_28), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (n_27), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (n_26), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (n_25), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (n_24), .A1 (hfn_ipo_n6), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (n_23), .A1 (hfn_ipo_n6), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (n_22), .A1 (hfn_ipo_n6), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (n_21), .A1 (hfn_ipo_n6), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (n_20), .A1 (hfn_ipo_n6), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (n_19), .A1 (hfn_ipo_n6), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (n_18), .A1 (hfn_ipo_n6), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (n_17), .A1 (hfn_ipo_n6), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (n_16), .A1 (hfn_ipo_n6), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (n_15), .A1 (hfn_ipo_n6), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (n_14), .A1 (hfn_ipo_n6), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (n_13), .A1 (hfn_ipo_n6), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (n_12), .A1 (hfn_ipo_n6), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (n_11), .A1 (hfn_ipo_n6), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (n_10), .A1 (hfn_ipo_n6), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (n_9), .A1 (hfn_ipo_n6), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (hfn_ipo_n6), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (hfn_ipo_n6), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (hfn_ipo_n6), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (hfn_ipo_n6), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (hfn_ipo_n6), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (hfn_ipo_n6), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (hfn_ipo_n6), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid0_10), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid0_10), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid0_10), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid0_10), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid0_10), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid0_10), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid0_10), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid0_10), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid0_10), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid0_10), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid0_10), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid0_10), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid0_10), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid0_10), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid0_10), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid0_10), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid0_10), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid0_10), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid0_10), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid0_10), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid0_10), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid0_10), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid0_10), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid0_10), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid0_10), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid0_10), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid0_10), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid0_10), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid0_10), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid0_10), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid0_10), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (out[31]), .CK (CTS_n_tid0_10), .D (n_33));
DFF_X1 \out_reg[32]  (.Q (out[32]), .CK (CTS_n_tid0_10), .D (n_34));
DFF_X1 \out_reg[33]  (.Q (out[33]), .CK (CTS_n_tid0_10), .D (n_35));
DFF_X1 \out_reg[34]  (.Q (out[34]), .CK (CTS_n_tid0_10), .D (n_36));
DFF_X1 \out_reg[35]  (.Q (out[35]), .CK (CTS_n_tid0_10), .D (n_37));
DFF_X1 \out_reg[36]  (.Q (out[36]), .CK (CTS_n_tid0_10), .D (n_38));
DFF_X1 \out_reg[37]  (.Q (out[37]), .CK (CTS_n_tid0_10), .D (n_39));
DFF_X1 \out_reg[38]  (.Q (out[38]), .CK (CTS_n_tid0_10), .D (n_40));
DFF_X1 \out_reg[39]  (.Q (out[39]), .CK (CTS_n_tid0_10), .D (n_41));
DFF_X1 \out_reg[40]  (.Q (out[40]), .CK (CTS_n_tid0_10), .D (n_42));
DFF_X1 \out_reg[41]  (.Q (out[41]), .CK (CTS_n_tid0_10), .D (n_43));
DFF_X1 \out_reg[42]  (.Q (out[42]), .CK (CTS_n_tid0_10), .D (n_44));
DFF_X1 \out_reg[43]  (.Q (out[43]), .CK (CTS_n_tid0_10), .D (n_45));
DFF_X1 \out_reg[44]  (.Q (out[44]), .CK (CTS_n_tid0_10), .D (n_46));
DFF_X1 \out_reg[45]  (.Q (out[45]), .CK (CTS_n_tid0_10), .D (n_47));
DFF_X1 \out_reg[46]  (.Q (out[46]), .CK (CTS_n_tid0_10), .D (n_48));
DFF_X1 \out_reg[47]  (.Q (out[47]), .CK (CTS_n_tid0_10), .D (n_49));
DFF_X1 \out_reg[48]  (.Q (out[48]), .CK (CTS_n_tid0_10), .D (n_50));
DFF_X1 \out_reg[49]  (.Q (out[49]), .CK (CTS_n_tid0_10), .D (n_51));
DFF_X1 \out_reg[50]  (.Q (out[50]), .CK (CTS_n_tid0_10), .D (n_52));
DFF_X1 \out_reg[51]  (.Q (out[51]), .CK (CTS_n_tid0_10), .D (n_53));
DFF_X1 \out_reg[52]  (.Q (out[52]), .CK (CTS_n_tid0_10), .D (n_54));
DFF_X1 \out_reg[53]  (.Q (out[53]), .CK (CTS_n_tid0_10), .D (n_55));
DFF_X1 \out_reg[54]  (.Q (out[54]), .CK (CTS_n_tid0_10), .D (n_56));
DFF_X1 \out_reg[55]  (.Q (out[55]), .CK (CTS_n_tid0_10), .D (n_57));
DFF_X1 \out_reg[56]  (.Q (out[56]), .CK (CTS_n_tid0_10), .D (n_58));
DFF_X1 \out_reg[57]  (.Q (out[57]), .CK (CTS_n_tid0_10), .D (n_59));
DFF_X1 \out_reg[58]  (.Q (out[58]), .CK (CTS_n_tid0_10), .D (n_60));
DFF_X1 \out_reg[59]  (.Q (out[59]), .CK (CTS_n_tid0_10), .D (n_61));
DFF_X1 \out_reg[60]  (.Q (out[60]), .CK (CTS_n_tid0_10), .D (n_62));
DFF_X1 \out_reg[61]  (.Q (out[61]), .CK (CTS_n_tid0_10), .D (n_63));
DFF_X1 \out_reg[62]  (.Q (out[62]), .CK (CTS_n_tid0_10), .D (n_64));
DFF_X1 \out_reg[63]  (.Q (out[63]), .CK (CTS_n_tid0_10), .D (n_65));
CLKGATE_X8 clk_gate_out_reg (.GCK (CTS_n_tid0_11), .CK (clk_CTS_1_PP_0), .E (n_1));
CLKBUF_X3 CTS_L3_c_tid0_11 (.Z (CTS_n_tid0_10), .A (CTS_n_tid0_11));
CLKBUF_X3 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_0_0));

endmodule //registerNbits__parameterized0

module datapath__0_26 (p_0, i_in2);

output [31:0] p_0;
input [31:0] i_in2;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (i_in2[25]));
INV_X1 i_63 (.ZN (n_32), .A (i_in2[21]));
INV_X1 i_62 (.ZN (n_31), .A (i_in2[14]));
INV_X1 i_61 (.ZN (n_30), .A (i_in2[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (i_in2[2]), .A2 (i_in2[1]), .A3 (i_in2[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (i_in2[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (i_in2[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (i_in2[5]), .A3 (i_in2[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (i_in2[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (i_in2[8]), .A3 (i_in2[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (i_in2[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (i_in2[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (i_in2[12]), .A3 (i_in2[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (i_in2[15]), .A3 (i_in2[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (i_in2[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (i_in2[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (i_in2[18]), .A3 (i_in2[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (i_in2[18]), .A3 (i_in2[19]), .A4 (i_in2[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (i_in2[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (i_in2[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (i_in2[23]), .A3 (i_in2[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (i_in2[26]), .A3 (i_in2[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (i_in2[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (i_in2[28]), .A3 (i_in2[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (i_in2[28]), .A3 (i_in2[29]), .A4 (i_in2[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (i_in2[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (i_in2[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (i_in2[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (i_in2[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (i_in2[27]), .B1 (n_9), .B2 (i_in2[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (i_in2[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (i_in2[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (i_in2[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (i_in2[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (i_in2[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (i_in2[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (i_in2[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (i_in2[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (i_in2[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (i_in2[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (i_in2[16]), .B1 (n_19), .B2 (i_in2[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (i_in2[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (i_in2[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (i_in2[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (i_in2[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (i_in2[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (i_in2[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (i_in2[9]), .B1 (n_25), .B2 (i_in2[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (i_in2[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (i_in2[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (i_in2[6]), .B1 (n_27), .B2 (i_in2[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (i_in2[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (i_in2[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (i_in2[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (i_in2[2]), .B1 (i_in2[1]), .B2 (i_in2[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (i_in2[1]), .B (i_in2[0]));

endmodule //datapath__0_26

module datapath__0_24 (p_0, i_in1);

output [31:0] p_0;
input [31:0] i_in1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (i_in1[25]));
INV_X1 i_63 (.ZN (n_32), .A (i_in1[21]));
INV_X1 i_62 (.ZN (n_31), .A (i_in1[14]));
INV_X1 i_61 (.ZN (n_30), .A (i_in1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (i_in1[2]), .A2 (i_in1[1]), .A3 (i_in1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (i_in1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (i_in1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (i_in1[5]), .A3 (i_in1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (i_in1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (i_in1[8]), .A3 (i_in1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (i_in1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (i_in1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (i_in1[12]), .A3 (i_in1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (i_in1[15]), .A3 (i_in1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (i_in1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (i_in1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (i_in1[18]), .A3 (i_in1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (i_in1[18]), .A3 (i_in1[19]), .A4 (i_in1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (i_in1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (i_in1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (i_in1[23]), .A3 (i_in1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (i_in1[26]), .A3 (i_in1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (i_in1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (i_in1[28]), .A3 (i_in1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (i_in1[28]), .A3 (i_in1[29]), .A4 (i_in1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (i_in1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (i_in1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (i_in1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (i_in1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (i_in1[27]), .B1 (n_9), .B2 (i_in1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (i_in1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (i_in1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (i_in1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (i_in1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (i_in1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (i_in1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (i_in1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (i_in1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (i_in1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (i_in1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (i_in1[16]), .B1 (n_19), .B2 (i_in1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (i_in1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (i_in1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (i_in1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (i_in1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (i_in1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (i_in1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (i_in1[9]), .B1 (n_25), .B2 (i_in1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (i_in1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (i_in1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (i_in1[6]), .B1 (n_27), .B2 (i_in1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (i_in1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (i_in1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (i_in1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (i_in1[2]), .B1 (i_in1[1]), .B2 (i_in1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (i_in1[1]), .B (i_in1[0]));

endmodule //datapath__0_24

module datapath__0_21 (p_0, out);

output [63:0] p_0;
input [63:0] out;
wire n_61;
wire n_0;
wire n_60;
wire n_59;
wire n_58;
wire n_1;
wire n_57;
wire n_56;
wire n_2;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_3;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_4;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_5;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;


INV_X1 i_135 (.ZN (n_72), .A (out[60]));
INV_X1 i_134 (.ZN (n_71), .A (out[55]));
INV_X1 i_133 (.ZN (n_70), .A (out[51]));
INV_X1 i_132 (.ZN (n_69), .A (out[42]));
INV_X1 i_131 (.ZN (n_68), .A (out[40]));
INV_X1 i_130 (.ZN (n_67), .A (out[36]));
INV_X1 i_129 (.ZN (n_66), .A (out[31]));
INV_X1 i_128 (.ZN (n_65), .A (out[26]));
INV_X1 i_127 (.ZN (n_64), .A (out[21]));
INV_X1 i_126 (.ZN (n_63), .A (out[13]));
INV_X1 i_125 (.ZN (n_62), .A (out[11]));
OR3_X1 i_124 (.ZN (n_61), .A1 (out[2]), .A2 (out[1]), .A3 (out[0]));
OR2_X1 i_123 (.ZN (n_60), .A1 (n_61), .A2 (out[3]));
OR2_X1 i_122 (.ZN (n_59), .A1 (n_60), .A2 (out[4]));
OR3_X1 i_121 (.ZN (n_58), .A1 (n_59), .A2 (out[5]), .A3 (out[6]));
OR2_X1 i_120 (.ZN (n_57), .A1 (n_58), .A2 (out[7]));
OR3_X1 i_119 (.ZN (n_56), .A1 (n_57), .A2 (out[8]), .A3 (out[9]));
NOR2_X1 i_118 (.ZN (n_55), .A1 (n_56), .A2 (out[10]));
NAND2_X1 i_117 (.ZN (n_54), .A1 (n_55), .A2 (n_62));
NOR2_X1 i_116 (.ZN (n_53), .A1 (n_54), .A2 (out[12]));
NAND2_X1 i_115 (.ZN (n_52), .A1 (n_53), .A2 (n_63));
OR3_X1 i_114 (.ZN (n_51), .A1 (n_52), .A2 (out[14]), .A3 (out[15]));
OR2_X1 i_113 (.ZN (n_50), .A1 (n_51), .A2 (out[16]));
OR2_X1 i_112 (.ZN (n_49), .A1 (n_50), .A2 (out[17]));
NOR2_X1 i_111 (.ZN (n_48), .A1 (n_49), .A2 (out[18]));
NOR3_X1 i_110 (.ZN (n_47), .A1 (n_49), .A2 (out[18]), .A3 (out[19]));
NOR4_X1 i_109 (.ZN (n_46), .A1 (n_49), .A2 (out[18]), .A3 (out[19]), .A4 (out[20]));
NAND2_X1 i_108 (.ZN (n_45), .A1 (n_46), .A2 (n_64));
OR2_X1 i_107 (.ZN (n_44), .A1 (n_45), .A2 (out[22]));
NOR2_X1 i_106 (.ZN (n_43), .A1 (n_44), .A2 (out[23]));
NOR3_X1 i_105 (.ZN (n_42), .A1 (n_44), .A2 (out[23]), .A3 (out[24]));
NOR4_X1 i_104 (.ZN (n_41), .A1 (n_44), .A2 (out[23]), .A3 (out[24]), .A4 (out[25]));
NAND2_X1 i_103 (.ZN (n_40), .A1 (n_41), .A2 (n_65));
OR2_X1 i_102 (.ZN (n_39), .A1 (n_40), .A2 (out[27]));
NOR2_X1 i_101 (.ZN (n_38), .A1 (n_39), .A2 (out[28]));
NOR3_X1 i_100 (.ZN (n_37), .A1 (n_39), .A2 (out[28]), .A3 (out[29]));
NOR4_X1 i_99 (.ZN (n_36), .A1 (n_39), .A2 (out[28]), .A3 (out[29]), .A4 (out[30]));
NAND2_X1 i_98 (.ZN (n_35), .A1 (n_36), .A2 (n_66));
OR2_X1 i_97 (.ZN (n_34), .A1 (n_35), .A2 (out[32]));
NOR2_X1 i_96 (.ZN (n_33), .A1 (n_34), .A2 (out[33]));
NOR3_X1 i_95 (.ZN (n_32), .A1 (n_34), .A2 (out[33]), .A3 (out[34]));
NOR4_X1 i_94 (.ZN (n_31), .A1 (n_34), .A2 (out[33]), .A3 (out[34]), .A4 (out[35]));
NAND2_X1 i_93 (.ZN (n_30), .A1 (n_31), .A2 (n_67));
OR2_X1 i_92 (.ZN (n_29), .A1 (n_30), .A2 (out[37]));
NOR2_X1 i_91 (.ZN (n_28), .A1 (n_29), .A2 (out[38]));
NOR3_X1 i_90 (.ZN (n_27), .A1 (n_29), .A2 (out[38]), .A3 (out[39]));
NAND2_X1 i_89 (.ZN (n_26), .A1 (n_27), .A2 (n_68));
NOR2_X1 i_88 (.ZN (n_25), .A1 (n_26), .A2 (out[41]));
NAND2_X1 i_87 (.ZN (n_24), .A1 (n_25), .A2 (n_69));
OR3_X1 i_86 (.ZN (n_23), .A1 (n_24), .A2 (out[43]), .A3 (out[44]));
OR2_X1 i_85 (.ZN (n_22), .A1 (n_23), .A2 (out[45]));
OR2_X1 i_84 (.ZN (n_21), .A1 (n_22), .A2 (out[46]));
OR2_X1 i_83 (.ZN (n_20), .A1 (n_21), .A2 (out[47]));
NOR2_X1 i_82 (.ZN (n_19), .A1 (n_20), .A2 (out[48]));
NOR3_X1 i_81 (.ZN (n_18), .A1 (n_20), .A2 (out[48]), .A3 (out[49]));
NOR4_X1 i_80 (.ZN (n_17), .A1 (n_20), .A2 (out[48]), .A3 (out[49]), .A4 (out[50]));
NAND2_X1 i_79 (.ZN (n_16), .A1 (n_17), .A2 (n_70));
NOR2_X1 i_78 (.ZN (n_15), .A1 (n_16), .A2 (out[52]));
NOR3_X1 i_77 (.ZN (n_14), .A1 (n_16), .A2 (out[52]), .A3 (out[53]));
NOR4_X1 i_76 (.ZN (n_13), .A1 (n_16), .A2 (out[52]), .A3 (out[53]), .A4 (out[54]));
NAND2_X1 i_75 (.ZN (n_12), .A1 (n_13), .A2 (n_71));
OR3_X1 i_74 (.ZN (n_11), .A1 (n_12), .A2 (out[56]), .A3 (out[57]));
NOR2_X1 i_73 (.ZN (n_10), .A1 (n_11), .A2 (out[58]));
NOR3_X1 i_72 (.ZN (n_9), .A1 (n_11), .A2 (out[58]), .A3 (out[59]));
NAND2_X1 i_71 (.ZN (n_8), .A1 (n_9), .A2 (n_72));
NOR2_X1 i_70 (.ZN (n_7), .A1 (n_8), .A2 (out[61]));
NOR3_X1 i_69 (.ZN (n_6), .A1 (n_8), .A2 (out[61]), .A3 (out[62]));
XNOR2_X1 i_68 (.ZN (p_0[63]), .A (out[63]), .B (n_6));
XNOR2_X1 i_67 (.ZN (p_0[62]), .A (out[62]), .B (n_7));
XOR2_X1 i_66 (.Z (p_0[61]), .A (out[61]), .B (n_8));
XNOR2_X1 i_65 (.ZN (p_0[60]), .A (out[60]), .B (n_9));
XNOR2_X1 i_64 (.ZN (p_0[59]), .A (out[59]), .B (n_10));
XOR2_X1 i_63 (.Z (p_0[58]), .A (out[58]), .B (n_11));
OAI21_X1 i_62 (.ZN (n_5), .A (out[57]), .B1 (n_12), .B2 (out[56]));
AND2_X1 i_61 (.ZN (p_0[57]), .A1 (n_11), .A2 (n_5));
XOR2_X1 i_60 (.Z (p_0[56]), .A (out[56]), .B (n_12));
XNOR2_X1 i_59 (.ZN (p_0[55]), .A (out[55]), .B (n_13));
XNOR2_X1 i_58 (.ZN (p_0[54]), .A (out[54]), .B (n_14));
XNOR2_X1 i_57 (.ZN (p_0[53]), .A (out[53]), .B (n_15));
XOR2_X1 i_56 (.Z (p_0[52]), .A (out[52]), .B (n_16));
XNOR2_X1 i_55 (.ZN (p_0[51]), .A (out[51]), .B (n_17));
XNOR2_X1 i_54 (.ZN (p_0[50]), .A (out[50]), .B (n_18));
XNOR2_X1 i_53 (.ZN (p_0[49]), .A (out[49]), .B (n_19));
XOR2_X1 i_52 (.Z (p_0[48]), .A (out[48]), .B (n_20));
XOR2_X1 i_51 (.Z (p_0[47]), .A (out[47]), .B (n_21));
XOR2_X1 i_50 (.Z (p_0[46]), .A (out[46]), .B (n_22));
XOR2_X1 i_49 (.Z (p_0[45]), .A (out[45]), .B (n_23));
OAI21_X1 i_48 (.ZN (n_4), .A (out[44]), .B1 (n_24), .B2 (out[43]));
AND2_X1 i_47 (.ZN (p_0[44]), .A1 (n_23), .A2 (n_4));
XOR2_X1 i_46 (.Z (p_0[43]), .A (out[43]), .B (n_24));
XNOR2_X1 i_45 (.ZN (p_0[42]), .A (out[42]), .B (n_25));
XOR2_X1 i_44 (.Z (p_0[41]), .A (out[41]), .B (n_26));
XNOR2_X1 i_43 (.ZN (p_0[40]), .A (out[40]), .B (n_27));
XNOR2_X1 i_42 (.ZN (p_0[39]), .A (out[39]), .B (n_28));
XOR2_X1 i_41 (.Z (p_0[38]), .A (out[38]), .B (n_29));
XOR2_X1 i_40 (.Z (p_0[37]), .A (out[37]), .B (n_30));
XNOR2_X1 i_39 (.ZN (p_0[36]), .A (out[36]), .B (n_31));
XNOR2_X1 i_38 (.ZN (p_0[35]), .A (out[35]), .B (n_32));
XNOR2_X1 i_37 (.ZN (p_0[34]), .A (out[34]), .B (n_33));
XOR2_X1 i_36 (.Z (p_0[33]), .A (out[33]), .B (n_34));
XOR2_X1 i_35 (.Z (p_0[32]), .A (out[32]), .B (n_35));
XNOR2_X1 i_34 (.ZN (p_0[31]), .A (out[31]), .B (n_36));
XNOR2_X1 i_33 (.ZN (p_0[30]), .A (out[30]), .B (n_37));
XNOR2_X1 i_32 (.ZN (p_0[29]), .A (out[29]), .B (n_38));
XOR2_X1 i_31 (.Z (p_0[28]), .A (out[28]), .B (n_39));
XOR2_X1 i_30 (.Z (p_0[27]), .A (out[27]), .B (n_40));
XNOR2_X1 i_29 (.ZN (p_0[26]), .A (out[26]), .B (n_41));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (out[25]), .B (n_42));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (out[24]), .B (n_43));
XOR2_X1 i_26 (.Z (p_0[23]), .A (out[23]), .B (n_44));
XOR2_X1 i_25 (.Z (p_0[22]), .A (out[22]), .B (n_45));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (out[21]), .B (n_46));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (out[20]), .B (n_47));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (out[19]), .B (n_48));
XOR2_X1 i_21 (.Z (p_0[18]), .A (out[18]), .B (n_49));
XOR2_X1 i_20 (.Z (p_0[17]), .A (out[17]), .B (n_50));
XOR2_X1 i_19 (.Z (p_0[16]), .A (out[16]), .B (n_51));
OAI21_X1 i_18 (.ZN (n_3), .A (out[15]), .B1 (n_52), .B2 (out[14]));
AND2_X1 i_17 (.ZN (p_0[15]), .A1 (n_51), .A2 (n_3));
XOR2_X1 i_16 (.Z (p_0[14]), .A (out[14]), .B (n_52));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (out[13]), .B (n_53));
XOR2_X1 i_14 (.Z (p_0[12]), .A (out[12]), .B (n_54));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (out[11]), .B (n_55));
XOR2_X1 i_12 (.Z (p_0[10]), .A (out[10]), .B (n_56));
OAI21_X1 i_11 (.ZN (n_2), .A (out[9]), .B1 (n_57), .B2 (out[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_56), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (out[8]), .B (n_57));
XOR2_X1 i_8 (.Z (p_0[7]), .A (out[7]), .B (n_58));
OAI21_X1 i_7 (.ZN (n_1), .A (out[6]), .B1 (n_59), .B2 (out[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_58), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (out[5]), .B (n_59));
XOR2_X1 i_4 (.Z (p_0[4]), .A (out[4]), .B (n_60));
XOR2_X1 i_3 (.Z (p_0[3]), .A (out[3]), .B (n_61));
OAI21_X1 i_2 (.ZN (n_0), .A (out[2]), .B1 (out[1]), .B2 (out[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_61), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (out[1]), .B (out[0]));

endmodule //datapath__0_21

module shifter (i_clk_CTS_1_PP_0, i_clk_CTS_1_PP_1, i_clk, i_rst, i_load, i_add, 
    i_shift, i_out, i_sign, i_adder, Q, A, o_lsb, o_out);

output [31:0] A;
output o_lsb;
output [63:0] o_out;
input [31:0] Q;
input i_add;
input [32:0] i_adder;
input i_clk;
input i_load;
input i_out;
input i_rst;
input i_shift;
input i_sign;
input i_clk_CTS_1_PP_0;
input i_clk_CTS_1_PP_1;
wire add_temp;
wire n_0_0;
wire n_0_1;
wire n_0_2;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_99;
wire CTS_n_tid0_14;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_1;
wire n_65;
wire n_2;
wire n_64;
wire n_3;
wire n_63;
wire n_4;
wire n_62;
wire n_5;
wire n_61;
wire n_6;
wire n_60;
wire n_7;
wire n_59;
wire n_8;
wire n_58;
wire n_9;
wire n_57;
wire n_10;
wire n_56;
wire n_11;
wire n_55;
wire n_12;
wire n_54;
wire n_13;
wire n_53;
wire n_14;
wire n_52;
wire n_15;
wire n_51;
wire n_16;
wire n_50;
wire n_17;
wire n_49;
wire n_18;
wire n_48;
wire n_19;
wire n_47;
wire n_20;
wire n_46;
wire n_21;
wire n_45;
wire n_22;
wire n_44;
wire n_23;
wire n_43;
wire n_24;
wire n_42;
wire n_25;
wire n_41;
wire n_26;
wire n_40;
wire n_27;
wire n_39;
wire n_28;
wire n_38;
wire n_29;
wire n_37;
wire n_30;
wire n_36;
wire n_31;
wire n_35;
wire n_32;
wire n_33;
wire n_34;
wire hfn_ipo_n9;
wire hfn_ipo_n10;
wire drc_ipo_n12;
wire drc_ipo_n11;
wire CTS_n_tid0_15;


INV_X1 i_0_202 (.ZN (n_0_71), .A (i_rst));
INV_X1 i_0_201 (.ZN (n_0_70), .A (i_load));
INV_X1 i_0_200 (.ZN (n_0_69), .A (i_add));
NAND2_X1 i_0_199 (.ZN (n_0_68), .A1 (n_0_69), .A2 (i_shift));
NAND3_X1 i_0_198 (.ZN (n_99), .A1 (n_0_71), .A2 (n_0_70), .A3 (n_0_68));
NOR3_X1 i_0_197 (.ZN (n_0_67), .A1 (n_0_68), .A2 (i_load), .A3 (i_rst));
AND2_X4 i_0_196 (.ZN (n_0_66), .A1 (add_temp), .A2 (drc_ipo_n11));
AND2_X1 i_0_195 (.ZN (n_98), .A1 (i_adder[32]), .A2 (n_0_66));
NOR4_X1 i_0_194 (.ZN (n_0_65), .A1 (n_0_68), .A2 (add_temp), .A3 (i_load), .A4 (i_rst));
AOI22_X1 i_0_193 (.ZN (n_0_64), .A1 (i_adder[31]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[31]));
INV_X1 i_0_192 (.ZN (n_97), .A (n_0_64));
AOI22_X1 i_0_191 (.ZN (n_0_63), .A1 (i_adder[30]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[30]));
INV_X1 i_0_190 (.ZN (n_96), .A (n_0_63));
AOI22_X1 i_0_189 (.ZN (n_0_62), .A1 (i_adder[29]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[29]));
INV_X1 i_0_188 (.ZN (n_95), .A (n_0_62));
AOI22_X1 i_0_187 (.ZN (n_0_61), .A1 (i_adder[28]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[28]));
INV_X1 i_0_186 (.ZN (n_94), .A (n_0_61));
AOI22_X1 i_0_185 (.ZN (n_0_60), .A1 (i_adder[27]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[27]));
INV_X1 i_0_184 (.ZN (n_93), .A (n_0_60));
AOI22_X1 i_0_183 (.ZN (n_0_59), .A1 (i_adder[26]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[26]));
INV_X1 i_0_182 (.ZN (n_92), .A (n_0_59));
AOI22_X1 i_0_181 (.ZN (n_0_58), .A1 (i_adder[25]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[25]));
INV_X1 i_0_180 (.ZN (n_91), .A (n_0_58));
AOI22_X1 i_0_179 (.ZN (n_0_57), .A1 (i_adder[24]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[24]));
INV_X1 i_0_178 (.ZN (n_90), .A (n_0_57));
AOI22_X1 i_0_177 (.ZN (n_0_56), .A1 (i_adder[23]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[23]));
INV_X1 i_0_176 (.ZN (n_89), .A (n_0_56));
AOI22_X1 i_0_175 (.ZN (n_0_55), .A1 (i_adder[22]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[22]));
INV_X1 i_0_174 (.ZN (n_88), .A (n_0_55));
AOI22_X1 i_0_173 (.ZN (n_0_54), .A1 (i_adder[21]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[21]));
INV_X1 i_0_172 (.ZN (n_87), .A (n_0_54));
AOI22_X1 i_0_171 (.ZN (n_0_53), .A1 (i_adder[20]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[20]));
INV_X1 i_0_170 (.ZN (n_86), .A (n_0_53));
AOI22_X1 i_0_169 (.ZN (n_0_52), .A1 (i_adder[19]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[19]));
INV_X1 i_0_168 (.ZN (n_85), .A (n_0_52));
AOI22_X1 i_0_167 (.ZN (n_0_51), .A1 (i_adder[18]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[18]));
INV_X1 i_0_166 (.ZN (n_84), .A (n_0_51));
AOI22_X1 i_0_165 (.ZN (n_0_50), .A1 (i_adder[17]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[17]));
INV_X1 i_0_164 (.ZN (n_83), .A (n_0_50));
AOI22_X1 i_0_163 (.ZN (n_0_49), .A1 (i_adder[16]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[16]));
INV_X1 i_0_162 (.ZN (n_82), .A (n_0_49));
AOI22_X1 i_0_161 (.ZN (n_0_48), .A1 (i_adder[15]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[15]));
INV_X1 i_0_160 (.ZN (n_81), .A (n_0_48));
AOI22_X1 i_0_159 (.ZN (n_0_47), .A1 (i_adder[14]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[14]));
INV_X1 i_0_158 (.ZN (n_80), .A (n_0_47));
AOI22_X1 i_0_157 (.ZN (n_0_46), .A1 (i_adder[13]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[13]));
INV_X1 i_0_156 (.ZN (n_79), .A (n_0_46));
AOI22_X1 i_0_155 (.ZN (n_0_45), .A1 (i_adder[12]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[12]));
INV_X1 i_0_154 (.ZN (n_78), .A (n_0_45));
AOI22_X1 i_0_153 (.ZN (n_0_44), .A1 (i_adder[11]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[11]));
INV_X1 i_0_152 (.ZN (n_77), .A (n_0_44));
AOI22_X1 i_0_151 (.ZN (n_0_43), .A1 (i_adder[10]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[10]));
INV_X1 i_0_150 (.ZN (n_76), .A (n_0_43));
AOI22_X1 i_0_149 (.ZN (n_0_42), .A1 (i_adder[9]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[9]));
INV_X1 i_0_148 (.ZN (n_75), .A (n_0_42));
AOI22_X1 i_0_147 (.ZN (n_0_41), .A1 (i_adder[8]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[8]));
INV_X1 i_0_146 (.ZN (n_74), .A (n_0_41));
AOI22_X1 i_0_145 (.ZN (n_0_40), .A1 (i_adder[7]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[7]));
INV_X1 i_0_144 (.ZN (n_73), .A (n_0_40));
AOI22_X1 i_0_143 (.ZN (n_0_39), .A1 (i_adder[6]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[6]));
INV_X1 i_0_142 (.ZN (n_72), .A (n_0_39));
AOI22_X1 i_0_141 (.ZN (n_0_38), .A1 (i_adder[5]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[5]));
INV_X1 i_0_140 (.ZN (n_71), .A (n_0_38));
AOI22_X1 i_0_139 (.ZN (n_0_37), .A1 (i_adder[4]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[4]));
INV_X1 i_0_138 (.ZN (n_70), .A (n_0_37));
AOI22_X1 i_0_137 (.ZN (n_0_36), .A1 (i_adder[3]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[3]));
INV_X1 i_0_136 (.ZN (n_69), .A (n_0_36));
AOI22_X1 i_0_135 (.ZN (n_0_35), .A1 (i_adder[2]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[2]));
INV_X1 i_0_134 (.ZN (n_68), .A (n_0_35));
AOI22_X1 i_0_133 (.ZN (n_0_34), .A1 (i_adder[1]), .A2 (n_0_66), .B1 (drc_ipo_n12), .B2 (A[1]));
INV_X1 i_0_132 (.ZN (n_67), .A (n_0_34));
NOR2_X4 i_0_131 (.ZN (n_0_33), .A1 (n_0_70), .A2 (i_rst));
AOI222_X1 i_0_130 (.ZN (n_0_32), .A1 (i_adder[0]), .A2 (n_0_66), .B1 (drc_ipo_n12)
    , .B2 (A[0]), .C1 (Q[31]), .C2 (n_0_33));
INV_X1 i_0_129 (.ZN (n_66), .A (n_0_32));
AOI22_X1 i_0_128 (.ZN (n_0_31), .A1 (n_1), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[30]));
INV_X1 i_0_127 (.ZN (n_65), .A (n_0_31));
AOI22_X1 i_0_126 (.ZN (n_0_30), .A1 (n_2), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[29]));
INV_X1 i_0_125 (.ZN (n_64), .A (n_0_30));
AOI22_X1 i_0_124 (.ZN (n_0_29), .A1 (n_3), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[28]));
INV_X1 i_0_123 (.ZN (n_63), .A (n_0_29));
AOI22_X1 i_0_122 (.ZN (n_0_28), .A1 (n_4), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[27]));
INV_X1 i_0_121 (.ZN (n_62), .A (n_0_28));
AOI22_X1 i_0_120 (.ZN (n_0_27), .A1 (n_5), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[26]));
INV_X1 i_0_119 (.ZN (n_61), .A (n_0_27));
AOI22_X1 i_0_118 (.ZN (n_0_26), .A1 (n_6), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[25]));
INV_X1 i_0_117 (.ZN (n_60), .A (n_0_26));
AOI22_X1 i_0_116 (.ZN (n_0_25), .A1 (n_7), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[24]));
INV_X1 i_0_115 (.ZN (n_59), .A (n_0_25));
AOI22_X1 i_0_114 (.ZN (n_0_24), .A1 (n_8), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[23]));
INV_X1 i_0_113 (.ZN (n_58), .A (n_0_24));
AOI22_X1 i_0_112 (.ZN (n_0_23), .A1 (n_9), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[22]));
INV_X1 i_0_111 (.ZN (n_57), .A (n_0_23));
AOI22_X1 i_0_110 (.ZN (n_0_22), .A1 (n_10), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[21]));
INV_X1 i_0_109 (.ZN (n_56), .A (n_0_22));
AOI22_X1 i_0_108 (.ZN (n_0_21), .A1 (n_11), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[20]));
INV_X1 i_0_107 (.ZN (n_55), .A (n_0_21));
AOI22_X1 i_0_106 (.ZN (n_0_20), .A1 (n_12), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[19]));
INV_X1 i_0_105 (.ZN (n_54), .A (n_0_20));
AOI22_X1 i_0_104 (.ZN (n_0_19), .A1 (n_13), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[18]));
INV_X1 i_0_103 (.ZN (n_53), .A (n_0_19));
AOI22_X1 i_0_102 (.ZN (n_0_18), .A1 (n_14), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[17]));
INV_X1 i_0_101 (.ZN (n_52), .A (n_0_18));
AOI22_X1 i_0_100 (.ZN (n_0_17), .A1 (n_15), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[16]));
INV_X1 i_0_99 (.ZN (n_51), .A (n_0_17));
AOI22_X1 i_0_98 (.ZN (n_0_16), .A1 (n_16), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[15]));
INV_X1 i_0_97 (.ZN (n_50), .A (n_0_16));
AOI22_X1 i_0_96 (.ZN (n_0_15), .A1 (n_17), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[14]));
INV_X1 i_0_95 (.ZN (n_49), .A (n_0_15));
AOI22_X1 i_0_94 (.ZN (n_0_14), .A1 (n_18), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[13]));
INV_X1 i_0_93 (.ZN (n_48), .A (n_0_14));
AOI22_X1 i_0_92 (.ZN (n_0_13), .A1 (n_19), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[12]));
INV_X1 i_0_91 (.ZN (n_47), .A (n_0_13));
AOI22_X1 i_0_90 (.ZN (n_0_12), .A1 (n_20), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[11]));
INV_X1 i_0_89 (.ZN (n_46), .A (n_0_12));
AOI22_X1 i_0_88 (.ZN (n_0_11), .A1 (n_21), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[10]));
INV_X1 i_0_87 (.ZN (n_45), .A (n_0_11));
AOI22_X1 i_0_86 (.ZN (n_0_10), .A1 (n_22), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[9]));
INV_X1 i_0_85 (.ZN (n_44), .A (n_0_10));
AOI22_X1 i_0_84 (.ZN (n_0_9), .A1 (n_23), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[8]));
INV_X1 i_0_83 (.ZN (n_43), .A (n_0_9));
AOI22_X1 i_0_82 (.ZN (n_0_8), .A1 (n_24), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[7]));
INV_X1 i_0_81 (.ZN (n_42), .A (n_0_8));
AOI22_X1 i_0_80 (.ZN (n_0_7), .A1 (n_25), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[6]));
INV_X1 i_0_79 (.ZN (n_41), .A (n_0_7));
AOI22_X1 i_0_78 (.ZN (n_0_6), .A1 (n_26), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[5]));
INV_X1 i_0_77 (.ZN (n_40), .A (n_0_6));
AOI22_X1 i_0_76 (.ZN (n_0_5), .A1 (n_27), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[4]));
INV_X1 i_0_75 (.ZN (n_39), .A (n_0_5));
AOI22_X1 i_0_74 (.ZN (n_0_4), .A1 (n_28), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[3]));
INV_X1 i_0_73 (.ZN (n_38), .A (n_0_4));
AOI22_X1 i_0_72 (.ZN (n_0_3), .A1 (n_29), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[2]));
INV_X1 i_0_71 (.ZN (n_37), .A (n_0_3));
AOI22_X1 i_0_70 (.ZN (n_0_2), .A1 (n_30), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[1]));
INV_X1 i_0_69 (.ZN (n_36), .A (n_0_2));
AOI22_X1 i_0_68 (.ZN (n_0_1), .A1 (n_31), .A2 (drc_ipo_n11), .B1 (n_0_33), .B2 (Q[0]));
INV_X1 i_0_67 (.ZN (n_35), .A (n_0_1));
AOI21_X1 i_0_66 (.ZN (n_0_0), .A (i_add), .B1 (i_shift), .B2 (add_temp));
OAI21_X1 i_0_65 (.ZN (n_34), .A (n_0_71), .B1 (i_load), .B2 (n_0_0));
NOR2_X1 i_0_64 (.ZN (n_33), .A1 (n_0_69), .A2 (i_rst));
AND2_X1 i_0_63 (.ZN (o_out[63]), .A1 (A[31]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_62 (.ZN (o_out[62]), .A1 (A[30]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_61 (.ZN (o_out[61]), .A1 (A[29]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_60 (.ZN (o_out[60]), .A1 (A[28]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_59 (.ZN (o_out[59]), .A1 (A[27]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_58 (.ZN (o_out[58]), .A1 (A[26]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_57 (.ZN (o_out[57]), .A1 (A[25]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_56 (.ZN (o_out[56]), .A1 (A[24]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_55 (.ZN (o_out[55]), .A1 (A[23]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_54 (.ZN (o_out[54]), .A1 (A[22]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_53 (.ZN (o_out[53]), .A1 (A[21]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_52 (.ZN (o_out[52]), .A1 (A[20]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_51 (.ZN (o_out[51]), .A1 (A[19]), .A2 (hfn_ipo_n10));
AND2_X1 i_0_50 (.ZN (o_out[50]), .A1 (A[18]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_49 (.ZN (o_out[49]), .A1 (A[17]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_48 (.ZN (o_out[48]), .A1 (A[16]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_47 (.ZN (o_out[47]), .A1 (A[15]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_46 (.ZN (o_out[46]), .A1 (A[14]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_45 (.ZN (o_out[45]), .A1 (A[13]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_44 (.ZN (o_out[44]), .A1 (A[12]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_43 (.ZN (o_out[43]), .A1 (A[11]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_42 (.ZN (o_out[42]), .A1 (A[10]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_41 (.ZN (o_out[41]), .A1 (A[9]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_40 (.ZN (o_out[40]), .A1 (A[8]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_39 (.ZN (o_out[39]), .A1 (A[7]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_38 (.ZN (o_out[38]), .A1 (A[6]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_37 (.ZN (o_out[37]), .A1 (A[5]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_36 (.ZN (o_out[36]), .A1 (A[4]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_35 (.ZN (o_out[35]), .A1 (A[3]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_34 (.ZN (o_out[34]), .A1 (A[2]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_33 (.ZN (o_out[33]), .A1 (A[1]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_32 (.ZN (o_out[32]), .A1 (A[0]), .A2 (hfn_ipo_n9));
AND2_X1 i_0_31 (.ZN (o_out[31]), .A1 (n_1), .A2 (hfn_ipo_n9));
AND2_X1 i_0_30 (.ZN (o_out[30]), .A1 (n_2), .A2 (hfn_ipo_n9));
AND2_X1 i_0_29 (.ZN (o_out[29]), .A1 (n_3), .A2 (hfn_ipo_n9));
AND2_X1 i_0_28 (.ZN (o_out[28]), .A1 (n_4), .A2 (hfn_ipo_n9));
AND2_X1 i_0_27 (.ZN (o_out[27]), .A1 (n_5), .A2 (hfn_ipo_n9));
AND2_X1 i_0_26 (.ZN (o_out[26]), .A1 (n_6), .A2 (hfn_ipo_n9));
AND2_X1 i_0_25 (.ZN (o_out[25]), .A1 (n_7), .A2 (hfn_ipo_n9));
AND2_X1 i_0_24 (.ZN (o_out[24]), .A1 (n_8), .A2 (hfn_ipo_n9));
AND2_X1 i_0_23 (.ZN (o_out[23]), .A1 (n_9), .A2 (hfn_ipo_n9));
AND2_X1 i_0_22 (.ZN (o_out[22]), .A1 (n_10), .A2 (hfn_ipo_n9));
AND2_X1 i_0_21 (.ZN (o_out[21]), .A1 (n_11), .A2 (hfn_ipo_n9));
AND2_X1 i_0_20 (.ZN (o_out[20]), .A1 (n_12), .A2 (hfn_ipo_n10));
AND2_X1 i_0_19 (.ZN (o_out[19]), .A1 (n_13), .A2 (hfn_ipo_n10));
AND2_X1 i_0_18 (.ZN (o_out[18]), .A1 (n_14), .A2 (hfn_ipo_n10));
AND2_X1 i_0_17 (.ZN (o_out[17]), .A1 (n_15), .A2 (hfn_ipo_n10));
AND2_X1 i_0_16 (.ZN (o_out[16]), .A1 (n_16), .A2 (hfn_ipo_n10));
AND2_X1 i_0_15 (.ZN (o_out[15]), .A1 (n_17), .A2 (hfn_ipo_n10));
AND2_X1 i_0_14 (.ZN (o_out[14]), .A1 (n_18), .A2 (hfn_ipo_n10));
AND2_X1 i_0_13 (.ZN (o_out[13]), .A1 (n_19), .A2 (hfn_ipo_n10));
AND2_X1 i_0_12 (.ZN (o_out[12]), .A1 (n_20), .A2 (hfn_ipo_n10));
AND2_X1 i_0_11 (.ZN (o_out[11]), .A1 (n_21), .A2 (hfn_ipo_n10));
AND2_X1 i_0_10 (.ZN (o_out[10]), .A1 (n_22), .A2 (hfn_ipo_n10));
AND2_X1 i_0_9 (.ZN (o_out[9]), .A1 (n_23), .A2 (hfn_ipo_n10));
AND2_X1 i_0_8 (.ZN (o_out[8]), .A1 (n_24), .A2 (hfn_ipo_n10));
AND2_X1 i_0_7 (.ZN (o_out[7]), .A1 (n_25), .A2 (hfn_ipo_n10));
AND2_X1 i_0_6 (.ZN (o_out[6]), .A1 (n_26), .A2 (hfn_ipo_n10));
AND2_X1 i_0_5 (.ZN (o_out[5]), .A1 (n_27), .A2 (hfn_ipo_n10));
AND2_X1 i_0_4 (.ZN (o_out[4]), .A1 (n_28), .A2 (hfn_ipo_n10));
AND2_X1 i_0_3 (.ZN (o_out[3]), .A1 (n_29), .A2 (hfn_ipo_n10));
AND2_X1 i_0_2 (.ZN (o_out[2]), .A1 (n_30), .A2 (hfn_ipo_n10));
AND2_X1 i_0_1 (.ZN (o_out[1]), .A1 (n_31), .A2 (hfn_ipo_n9));
AND2_X1 i_0_0 (.ZN (o_out[0]), .A1 (o_lsb), .A2 (hfn_ipo_n9));
MUX2_X1 add_temp_reg_enable_mux_0 (.Z (n_32), .A (add_temp), .B (n_33), .S (n_34));
DFF_X1 add_temp_reg (.Q (add_temp), .CK (i_clk_CTS_1_PP_0), .D (n_32));
DFF_X1 \temp_reg[0]  (.Q (o_lsb), .CK (CTS_n_tid0_14), .D (n_35));
DFF_X1 \temp_reg[1]  (.Q (n_31), .CK (CTS_n_tid0_14), .D (n_36));
DFF_X1 \temp_reg[2]  (.Q (n_30), .CK (CTS_n_tid0_14), .D (n_37));
DFF_X1 \temp_reg[3]  (.Q (n_29), .CK (CTS_n_tid0_14), .D (n_38));
DFF_X1 \temp_reg[4]  (.Q (n_28), .CK (CTS_n_tid0_14), .D (n_39));
DFF_X1 \temp_reg[5]  (.Q (n_27), .CK (CTS_n_tid0_14), .D (n_40));
DFF_X1 \temp_reg[6]  (.Q (n_26), .CK (CTS_n_tid0_14), .D (n_41));
DFF_X1 \temp_reg[7]  (.Q (n_25), .CK (CTS_n_tid0_14), .D (n_42));
DFF_X1 \temp_reg[8]  (.Q (n_24), .CK (CTS_n_tid0_14), .D (n_43));
DFF_X1 \temp_reg[9]  (.Q (n_23), .CK (CTS_n_tid0_14), .D (n_44));
DFF_X1 \temp_reg[10]  (.Q (n_22), .CK (CTS_n_tid0_14), .D (n_45));
DFF_X1 \temp_reg[11]  (.Q (n_21), .CK (CTS_n_tid0_14), .D (n_46));
DFF_X1 \temp_reg[12]  (.Q (n_20), .CK (CTS_n_tid0_14), .D (n_47));
DFF_X1 \temp_reg[13]  (.Q (n_19), .CK (CTS_n_tid0_14), .D (n_48));
DFF_X1 \temp_reg[14]  (.Q (n_18), .CK (CTS_n_tid0_14), .D (n_49));
DFF_X1 \temp_reg[15]  (.Q (n_17), .CK (CTS_n_tid0_14), .D (n_50));
DFF_X1 \temp_reg[16]  (.Q (n_16), .CK (CTS_n_tid0_14), .D (n_51));
DFF_X1 \temp_reg[17]  (.Q (n_15), .CK (CTS_n_tid0_14), .D (n_52));
DFF_X1 \temp_reg[18]  (.Q (n_14), .CK (CTS_n_tid0_14), .D (n_53));
DFF_X1 \temp_reg[19]  (.Q (n_13), .CK (CTS_n_tid0_14), .D (n_54));
DFF_X1 \temp_reg[20]  (.Q (n_12), .CK (CTS_n_tid0_14), .D (n_55));
DFF_X1 \temp_reg[21]  (.Q (n_11), .CK (CTS_n_tid0_14), .D (n_56));
DFF_X1 \temp_reg[22]  (.Q (n_10), .CK (CTS_n_tid0_14), .D (n_57));
DFF_X1 \temp_reg[23]  (.Q (n_9), .CK (CTS_n_tid0_14), .D (n_58));
DFF_X1 \temp_reg[24]  (.Q (n_8), .CK (CTS_n_tid0_14), .D (n_59));
DFF_X1 \temp_reg[25]  (.Q (n_7), .CK (CTS_n_tid0_14), .D (n_60));
DFF_X1 \temp_reg[26]  (.Q (n_6), .CK (CTS_n_tid0_14), .D (n_61));
DFF_X1 \temp_reg[27]  (.Q (n_5), .CK (CTS_n_tid0_14), .D (n_62));
DFF_X1 \temp_reg[28]  (.Q (n_4), .CK (CTS_n_tid0_14), .D (n_63));
DFF_X1 \temp_reg[29]  (.Q (n_3), .CK (CTS_n_tid0_14), .D (n_64));
DFF_X1 \temp_reg[30]  (.Q (n_2), .CK (CTS_n_tid0_14), .D (n_65));
DFF_X1 \temp_reg[31]  (.Q (n_1), .CK (CTS_n_tid0_14), .D (n_66));
DFF_X1 \temp_reg[32]  (.Q (A[0]), .CK (CTS_n_tid0_14), .D (n_67));
DFF_X1 \temp_reg[33]  (.Q (A[1]), .CK (CTS_n_tid0_14), .D (n_68));
DFF_X1 \temp_reg[34]  (.Q (A[2]), .CK (CTS_n_tid0_14), .D (n_69));
DFF_X1 \temp_reg[35]  (.Q (A[3]), .CK (CTS_n_tid0_14), .D (n_70));
DFF_X1 \temp_reg[36]  (.Q (A[4]), .CK (CTS_n_tid0_14), .D (n_71));
DFF_X1 \temp_reg[37]  (.Q (A[5]), .CK (CTS_n_tid0_14), .D (n_72));
DFF_X1 \temp_reg[38]  (.Q (A[6]), .CK (CTS_n_tid0_14), .D (n_73));
DFF_X1 \temp_reg[39]  (.Q (A[7]), .CK (CTS_n_tid0_14), .D (n_74));
DFF_X1 \temp_reg[40]  (.Q (A[8]), .CK (CTS_n_tid0_14), .D (n_75));
DFF_X1 \temp_reg[41]  (.Q (A[9]), .CK (CTS_n_tid0_14), .D (n_76));
DFF_X1 \temp_reg[42]  (.Q (A[10]), .CK (CTS_n_tid0_14), .D (n_77));
DFF_X1 \temp_reg[43]  (.Q (A[11]), .CK (CTS_n_tid0_14), .D (n_78));
DFF_X1 \temp_reg[44]  (.Q (A[12]), .CK (CTS_n_tid0_14), .D (n_79));
DFF_X1 \temp_reg[45]  (.Q (A[13]), .CK (CTS_n_tid0_14), .D (n_80));
DFF_X1 \temp_reg[46]  (.Q (A[14]), .CK (CTS_n_tid0_14), .D (n_81));
DFF_X1 \temp_reg[47]  (.Q (A[15]), .CK (CTS_n_tid0_14), .D (n_82));
DFF_X1 \temp_reg[48]  (.Q (A[16]), .CK (CTS_n_tid0_14), .D (n_83));
DFF_X1 \temp_reg[49]  (.Q (A[17]), .CK (CTS_n_tid0_14), .D (n_84));
DFF_X1 \temp_reg[50]  (.Q (A[18]), .CK (CTS_n_tid0_14), .D (n_85));
DFF_X1 \temp_reg[51]  (.Q (A[19]), .CK (CTS_n_tid0_14), .D (n_86));
DFF_X1 \temp_reg[52]  (.Q (A[20]), .CK (CTS_n_tid0_14), .D (n_87));
DFF_X1 \temp_reg[53]  (.Q (A[21]), .CK (CTS_n_tid0_14), .D (n_88));
DFF_X1 \temp_reg[54]  (.Q (A[22]), .CK (CTS_n_tid0_14), .D (n_89));
DFF_X1 \temp_reg[55]  (.Q (A[23]), .CK (CTS_n_tid0_14), .D (n_90));
DFF_X1 \temp_reg[56]  (.Q (A[24]), .CK (CTS_n_tid0_14), .D (n_91));
DFF_X1 \temp_reg[57]  (.Q (A[25]), .CK (CTS_n_tid0_14), .D (n_92));
DFF_X1 \temp_reg[58]  (.Q (A[26]), .CK (CTS_n_tid0_14), .D (n_93));
DFF_X1 \temp_reg[59]  (.Q (A[27]), .CK (CTS_n_tid0_14), .D (n_94));
DFF_X1 \temp_reg[60]  (.Q (A[28]), .CK (CTS_n_tid0_14), .D (n_95));
DFF_X1 \temp_reg[61]  (.Q (A[29]), .CK (CTS_n_tid0_14), .D (n_96));
DFF_X1 \temp_reg[62]  (.Q (A[30]), .CK (CTS_n_tid0_14), .D (n_97));
DFF_X1 \temp_reg[63]  (.Q (A[31]), .CK (CTS_n_tid0_14), .D (n_98));
CLKGATE_X8 clk_gate_temp_reg (.GCK (CTS_n_tid0_15), .CK (i_clk_CTS_1_PP_1), .E (n_99));
CLKBUF_X1 hfn_ipo_c9 (.Z (hfn_ipo_n9), .A (i_out));
CLKBUF_X1 hfn_ipo_c10 (.Z (hfn_ipo_n10), .A (i_out));
CLKBUF_X2 drc_ipo_c12 (.Z (drc_ipo_n12), .A (n_0_65));
BUF_X4 drc_ipo_c11 (.Z (drc_ipo_n11), .A (n_0_67));
CLKBUF_X3 CTS_L3_c_tid0_15 (.Z (CTS_n_tid0_14), .A (CTS_n_tid0_15));

endmodule //shifter

module datapath (i_in2, i_in1, o_out1);

output [32:0] o_out1;
input [31:0] i_in1;
input [31:0] i_in2;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;


FA_X1 i_31 (.CO (o_out1[32]), .S (o_out1[31]), .A (i_in2[31]), .B (i_in1[31]), .CI (n_30));
FA_X1 i_30 (.CO (n_30), .S (o_out1[30]), .A (i_in2[30]), .B (i_in1[30]), .CI (n_29));
FA_X1 i_29 (.CO (n_29), .S (o_out1[29]), .A (i_in2[29]), .B (i_in1[29]), .CI (n_28));
FA_X1 i_28 (.CO (n_28), .S (o_out1[28]), .A (i_in2[28]), .B (i_in1[28]), .CI (n_27));
FA_X1 i_27 (.CO (n_27), .S (o_out1[27]), .A (i_in2[27]), .B (i_in1[27]), .CI (n_26));
FA_X1 i_26 (.CO (n_26), .S (o_out1[26]), .A (i_in2[26]), .B (i_in1[26]), .CI (n_25));
FA_X1 i_25 (.CO (n_25), .S (o_out1[25]), .A (i_in2[25]), .B (i_in1[25]), .CI (n_24));
FA_X1 i_24 (.CO (n_24), .S (o_out1[24]), .A (i_in2[24]), .B (i_in1[24]), .CI (n_23));
FA_X1 i_23 (.CO (n_23), .S (o_out1[23]), .A (i_in2[23]), .B (i_in1[23]), .CI (n_22));
FA_X1 i_22 (.CO (n_22), .S (o_out1[22]), .A (i_in2[22]), .B (i_in1[22]), .CI (n_21));
FA_X1 i_21 (.CO (n_21), .S (o_out1[21]), .A (i_in2[21]), .B (i_in1[21]), .CI (n_20));
FA_X1 i_20 (.CO (n_20), .S (o_out1[20]), .A (i_in2[20]), .B (i_in1[20]), .CI (n_19));
FA_X1 i_19 (.CO (n_19), .S (o_out1[19]), .A (i_in2[19]), .B (i_in1[19]), .CI (n_18));
FA_X1 i_18 (.CO (n_18), .S (o_out1[18]), .A (i_in2[18]), .B (i_in1[18]), .CI (n_17));
FA_X1 i_17 (.CO (n_17), .S (o_out1[17]), .A (i_in2[17]), .B (i_in1[17]), .CI (n_16));
FA_X1 i_16 (.CO (n_16), .S (o_out1[16]), .A (i_in2[16]), .B (i_in1[16]), .CI (n_15));
FA_X1 i_15 (.CO (n_15), .S (o_out1[15]), .A (i_in2[15]), .B (i_in1[15]), .CI (n_14));
FA_X1 i_14 (.CO (n_14), .S (o_out1[14]), .A (i_in2[14]), .B (i_in1[14]), .CI (n_13));
FA_X1 i_13 (.CO (n_13), .S (o_out1[13]), .A (i_in2[13]), .B (i_in1[13]), .CI (n_12));
FA_X1 i_12 (.CO (n_12), .S (o_out1[12]), .A (i_in2[12]), .B (i_in1[12]), .CI (n_11));
FA_X1 i_11 (.CO (n_11), .S (o_out1[11]), .A (i_in2[11]), .B (i_in1[11]), .CI (n_10));
FA_X1 i_10 (.CO (n_10), .S (o_out1[10]), .A (i_in2[10]), .B (i_in1[10]), .CI (n_9));
FA_X1 i_9 (.CO (n_9), .S (o_out1[9]), .A (i_in2[9]), .B (i_in1[9]), .CI (n_8));
FA_X1 i_8 (.CO (n_8), .S (o_out1[8]), .A (i_in2[8]), .B (i_in1[8]), .CI (n_7));
FA_X1 i_7 (.CO (n_7), .S (o_out1[7]), .A (i_in2[7]), .B (i_in1[7]), .CI (n_6));
FA_X1 i_6 (.CO (n_6), .S (o_out1[6]), .A (i_in2[6]), .B (i_in1[6]), .CI (n_5));
FA_X1 i_5 (.CO (n_5), .S (o_out1[5]), .A (i_in2[5]), .B (i_in1[5]), .CI (n_4));
FA_X1 i_4 (.CO (n_4), .S (o_out1[4]), .A (i_in2[4]), .B (i_in1[4]), .CI (n_3));
FA_X1 i_3 (.CO (n_3), .S (o_out1[3]), .A (i_in2[3]), .B (i_in1[3]), .CI (n_2));
FA_X1 i_2 (.CO (n_2), .S (o_out1[2]), .A (i_in2[2]), .B (i_in1[2]), .CI (n_1));
FA_X1 i_1 (.CO (n_1), .S (o_out1[1]), .A (i_in2[1]), .B (i_in1[1]), .CI (n_0));
HA_X1 i_0 (.CO (n_0), .S (o_out1[0]), .A (i_in2[0]), .B (i_in1[0]));

endmodule //datapath

module adder (i_in1, i_in2, o_out1);

output [32:0] o_out1;
input [31:0] i_in1;
input [31:0] i_in2;


datapath i_0 (.o_out1 ({o_out1[32], o_out1[31], o_out1[30], o_out1[29], o_out1[28], 
    o_out1[27], o_out1[26], o_out1[25], o_out1[24], o_out1[23], o_out1[22], o_out1[21], 
    o_out1[20], o_out1[19], o_out1[18], o_out1[17], o_out1[16], o_out1[15], o_out1[14], 
    o_out1[13], o_out1[12], o_out1[11], o_out1[10], o_out1[9], o_out1[8], o_out1[7], 
    o_out1[6], o_out1[5], o_out1[4], o_out1[3], o_out1[2], o_out1[1], o_out1[0]})
    , .i_in1 ({i_in1[31], i_in1[30], i_in1[29], i_in1[28], i_in1[27], i_in1[26], 
    i_in1[25], i_in1[24], i_in1[23], i_in1[22], i_in1[21], i_in1[20], i_in1[19], 
    i_in1[18], i_in1[17], i_in1[16], i_in1[15], i_in1[14], i_in1[13], i_in1[12], 
    i_in1[11], i_in1[10], i_in1[9], i_in1[8], i_in1[7], i_in1[6], i_in1[5], i_in1[4], 
    i_in1[3], i_in1[2], i_in1[1], i_in1[0]}), .i_in2 ({i_in2[31], i_in2[30], i_in2[29], 
    i_in2[28], i_in2[27], i_in2[26], i_in2[25], i_in2[24], i_in2[23], i_in2[22], 
    i_in2[21], i_in2[20], i_in2[19], i_in2[18], i_in2[17], i_in2[16], i_in2[15], 
    i_in2[14], i_in2[13], i_in2[12], i_in2[11], i_in2[10], i_in2[9], i_in2[8], i_in2[7], 
    i_in2[6], i_in2[5], i_in2[4], i_in2[3], i_in2[2], i_in2[1], i_in2[0]}));

endmodule //adder

module controller (i_clk_CTS_1_PP_0, i_clk_CTS_1_PP_1, i_clk, i_rst, i_lsb, o_load, 
    o_add, o_shift, o_out);

output o_add;
output o_load;
output o_out;
output o_shift;
output i_clk_CTS_1_PP_0;
input i_clk;
input i_lsb;
input i_rst;
input i_clk_CTS_1_PP_1;
wire start;
wire \state[2] ;
wire \state[1] ;
wire \state[0] ;
wire n_0_3;
wire n_0_0;
wire n_0_4;
wire n_0_1;
wire n_0_5;
wire n_0_2;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_24;
wire n_1;
wire n_23;
wire n_21;
wire n_20;
wire n_0;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_19;
wire n_18;
wire n_13;
wire n_2;
wire n_12;
wire n_3;
wire n_11;
wire n_4;
wire n_10;
wire n_5;
wire n_9;
wire n_6;
wire n_8;
wire n_7;
wire n_22;


INV_X1 i_0_34 (.ZN (n_0_22), .A (i_rst));
INV_X1 i_0_33 (.ZN (n_0_21), .A (\state[0] ));
INV_X1 i_0_32 (.ZN (n_0_20), .A (i_lsb));
INV_X1 i_0_31 (.ZN (n_0_19), .A (start));
NOR2_X1 i_0_30 (.ZN (n_0_18), .A1 (i_rst), .A2 (\state[2] ));
INV_X1 i_0_29 (.ZN (n_0_17), .A (n_0_18));
OR2_X1 i_0_28 (.ZN (n_0_16), .A1 (\state[1] ), .A2 (\state[0] ));
NOR3_X1 i_0_27 (.ZN (n_24), .A1 (n_0_17), .A2 (n_0_16), .A3 (start));
NAND2_X1 i_0_26 (.ZN (n_0_15), .A1 (n_0_22), .A2 (\state[2] ));
INV_X1 i_0_25 (.ZN (n_23), .A (n_0_15));
NAND2_X1 i_0_24 (.ZN (n_22), .A1 (n_0_16), .A2 (n_23));
NAND2_X1 i_0_23 (.ZN (n_0_14), .A1 (\state[1] ), .A2 (n_0_18));
NOR2_X1 i_0_22 (.ZN (n_21), .A1 (n_0_21), .A2 (n_0_14));
NOR3_X1 i_0_21 (.ZN (n_20), .A1 (\state[1] ), .A2 (n_0_21), .A3 (n_0_17));
AOI21_X1 i_0_20 (.ZN (n_0_13), .A (i_rst), .B1 (n_2), .B2 (\state[2] ));
INV_X1 i_0_19 (.ZN (n_0_12), .A (n_0_13));
AOI21_X1 i_0_18 (.ZN (n_19), .A (n_0_18), .B1 (n_0_22), .B2 (n_0_16));
AOI21_X1 i_0_17 (.ZN (n_17), .A (n_0_13), .B1 (n_0_22), .B2 (n_0_16));
OAI21_X1 i_0_16 (.ZN (n_0_11), .A (\state[1] ), .B1 (\state[0] ), .B2 (n_0_20));
NOR2_X1 i_0_15 (.ZN (n_16), .A1 (n_0_17), .A2 (n_0_11));
AOI21_X1 i_0_14 (.ZN (n_0_10), .A (\state[2] ), .B1 (n_0_16), .B2 (n_0_11));
NOR2_X1 i_0_13 (.ZN (n_15), .A1 (n_0_12), .A2 (n_0_10));
OAI33_X1 i_0_12 (.ZN (n_14), .A1 (n_0_19), .A2 (n_0_17), .A3 (n_0_16), .B1 (\state[0] )
    , .B2 (n_0_20), .B3 (n_0_14));
NOR3_X1 i_0_11 (.ZN (n_0_9), .A1 (n_2), .A2 (n_0_16), .A3 (n_0_15));
INV_X1 i_0_10 (.ZN (n_0_8), .A (n_0_9));
AND2_X1 i_0_9 (.ZN (n_13), .A1 (n_0_7), .A2 (n_0_9));
AND2_X1 i_0_8 (.ZN (n_12), .A1 (n_0_6), .A2 (n_0_9));
AND2_X1 i_0_7 (.ZN (n_11), .A1 (n_0_5), .A2 (n_0_9));
AND2_X1 i_0_6 (.ZN (n_10), .A1 (n_0_4), .A2 (n_0_9));
AND2_X1 i_0_5 (.ZN (n_9), .A1 (n_0_3), .A2 (n_0_9));
NOR2_X1 i_0_4 (.ZN (n_8), .A1 (n_7), .A2 (n_0_8));
HA_X1 i_0_3 (.CO (n_0_7), .S (n_0_6), .A (n_3), .B (n_0_2));
HA_X1 i_0_2 (.CO (n_0_2), .S (n_0_5), .A (n_4), .B (n_0_1));
HA_X1 i_0_1 (.CO (n_0_1), .S (n_0_4), .A (n_5), .B (n_0_0));
HA_X1 i_0_0 (.CO (n_0_0), .S (n_0_3), .A (n_6), .B (n_7));
CLKGATE_X1 clk_gate_o_out_reg (.GCK (n_1), .CK (i_clk_CTS_1_PP_1), .E (n_22));
DFF_X1 \count_reg[0]  (.Q (n_7), .CK (n_18), .D (n_8));
DFF_X1 \count_reg[1]  (.Q (n_6), .CK (n_18), .D (n_9));
DFF_X1 \count_reg[2]  (.Q (n_5), .CK (n_18), .D (n_10));
DFF_X1 \count_reg[3]  (.Q (n_4), .CK (n_18), .D (n_11));
DFF_X1 \count_reg[4]  (.Q (n_3), .CK (n_18), .D (n_12));
DFF_X1 \count_reg[5]  (.Q (n_2), .CK (n_18), .D (n_13));
CLKGATE_X1 clk_gate_count_reg (.GCK (n_18), .CK (i_clk_CTS_1_PP_0), .E (n_19));
DFF_X1 \state_reg[0]  (.Q (\state[0] ), .CK (n_1), .D (n_14));
DFF_X1 \state_reg[1]  (.Q (\state[1] ), .CK (n_1), .D (n_15));
DFF_X1 \state_reg[2]  (.Q (\state[2] ), .CK (n_1), .D (n_16));
MUX2_X1 start_reg_enable_mux_0 (.Z (n_0), .A (start), .B (i_rst), .S (n_17));
DFF_X1 start_reg (.Q (start), .CK (i_clk_CTS_1_PP_0), .D (n_0));
DFF_X1 o_load_reg (.Q (o_load), .CK (n_1), .D (n_20));
DFF_X1 o_add_reg (.Q (o_add), .CK (n_1), .D (n_21));
DFF_X1 o_shift_reg (.Q (o_shift), .CK (n_1), .D (n_23));
DFF_X1 o_out_reg (.Q (o_out), .CK (n_1), .D (n_24));
CLKBUF_X1 CTS_L3_c_tid1_12 (.Z (i_clk_CTS_1_PP_0), .A (i_clk_CTS_1_PP_1));

endmodule //controller

module multunit (i_clk_CTS_1_PP_0, i_clk_CTS_1_PP_2, i_clk, i_rst, i_in1, i_in2, 
    o_out1);

output [63:0] o_out1;
input i_clk;
input [31:0] i_in1;
input [31:0] i_in2;
input i_rst;
input i_clk_CTS_1_PP_0;
input i_clk_CTS_1_PP_2;
wire CTS_n_tid1_9;
wire out_ready;
wire shift;
wire add;
wire load;
wire \add_out[32] ;
wire \add_out[31] ;
wire \add_out[30] ;
wire \add_out[29] ;
wire \add_out[28] ;
wire \add_out[27] ;
wire \add_out[26] ;
wire \add_out[25] ;
wire \add_out[24] ;
wire \add_out[23] ;
wire \add_out[22] ;
wire \add_out[21] ;
wire \add_out[20] ;
wire \add_out[19] ;
wire \add_out[18] ;
wire \add_out[17] ;
wire \add_out[16] ;
wire \add_out[15] ;
wire \add_out[14] ;
wire \add_out[13] ;
wire \add_out[12] ;
wire \add_out[11] ;
wire \add_out[10] ;
wire \add_out[9] ;
wire \add_out[8] ;
wire \add_out[7] ;
wire \add_out[6] ;
wire \add_out[5] ;
wire \add_out[4] ;
wire \add_out[3] ;
wire \add_out[2] ;
wire \add_out[1] ;
wire \add_out[0] ;
wire \out[63] ;
wire \out[62] ;
wire \out[61] ;
wire \out[60] ;
wire \out[59] ;
wire \out[58] ;
wire \out[57] ;
wire \out[56] ;
wire \out[55] ;
wire \out[54] ;
wire \out[53] ;
wire \out[52] ;
wire \out[51] ;
wire \out[50] ;
wire \out[49] ;
wire \out[48] ;
wire \out[47] ;
wire \out[46] ;
wire \out[45] ;
wire \out[44] ;
wire \out[43] ;
wire \out[42] ;
wire \out[41] ;
wire \out[40] ;
wire \out[39] ;
wire \out[38] ;
wire \out[37] ;
wire \out[36] ;
wire \out[35] ;
wire \out[34] ;
wire \out[33] ;
wire \out[32] ;
wire \out[31] ;
wire \out[30] ;
wire \out[29] ;
wire \out[28] ;
wire \out[27] ;
wire \out[26] ;
wire \out[25] ;
wire \out[24] ;
wire \out[23] ;
wire \out[22] ;
wire \out[21] ;
wire \out[20] ;
wire \out[19] ;
wire \out[18] ;
wire \out[17] ;
wire \out[16] ;
wire \out[15] ;
wire \out[14] ;
wire \out[13] ;
wire \out[12] ;
wire \out[11] ;
wire \out[10] ;
wire \out[9] ;
wire \out[8] ;
wire \out[7] ;
wire \out[6] ;
wire \out[5] ;
wire \out[4] ;
wire \out[3] ;
wire \out[2] ;
wire \out[1] ;
wire lsb;
wire \A[31] ;
wire \A[30] ;
wire \A[29] ;
wire \A[28] ;
wire \A[27] ;
wire \A[26] ;
wire \A[25] ;
wire \A[24] ;
wire \A[23] ;
wire \A[22] ;
wire \A[21] ;
wire \A[20] ;
wire \A[19] ;
wire \A[18] ;
wire \A[17] ;
wire \A[16] ;
wire \A[15] ;
wire \A[14] ;
wire \A[13] ;
wire \A[12] ;
wire \A[11] ;
wire \A[10] ;
wire \A[9] ;
wire \A[8] ;
wire \A[7] ;
wire \A[6] ;
wire \A[5] ;
wire \A[4] ;
wire \A[3] ;
wire \A[2] ;
wire \A[1] ;
wire \A[0] ;
wire n_1_0;
wire \M[31] ;
wire \M[30] ;
wire \M[29] ;
wire \M[28] ;
wire \M[27] ;
wire \M[26] ;
wire \M[25] ;
wire \M[24] ;
wire \M[23] ;
wire \M[22] ;
wire \M[21] ;
wire \M[20] ;
wire \M[19] ;
wire \M[18] ;
wire \M[17] ;
wire \M[16] ;
wire \M[15] ;
wire \M[14] ;
wire \M[13] ;
wire \M[12] ;
wire \M[11] ;
wire \M[10] ;
wire \M[9] ;
wire \M[8] ;
wire \M[7] ;
wire \M[6] ;
wire \M[5] ;
wire \M[4] ;
wire \M[3] ;
wire \M[2] ;
wire \M[1] ;
wire hfn_ipo_n6;
wire \Q[31] ;
wire \Q[30] ;
wire \Q[29] ;
wire \Q[28] ;
wire \Q[27] ;
wire \Q[26] ;
wire \Q[25] ;
wire \Q[24] ;
wire \Q[23] ;
wire \Q[22] ;
wire \Q[21] ;
wire \Q[20] ;
wire \Q[19] ;
wire \Q[18] ;
wire \Q[17] ;
wire \Q[16] ;
wire \Q[15] ;
wire \Q[14] ;
wire \Q[13] ;
wire \Q[12] ;
wire \Q[11] ;
wire \Q[10] ;
wire \Q[9] ;
wire \Q[8] ;
wire \Q[7] ;
wire \Q[6] ;
wire \Q[5] ;
wire \Q[4] ;
wire \Q[3] ;
wire \Q[2] ;
wire \Q[1] ;
wire hfn_ipo_n5;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire n_1;
wire n_0;
wire uc_0;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire uc_1;
wire n_124;
wire n_123;
wire n_122;
wire n_121;
wire n_120;
wire n_119;
wire n_118;
wire n_117;
wire n_116;
wire n_115;
wire n_114;
wire n_113;
wire n_112;
wire n_111;
wire n_110;
wire n_109;
wire n_108;
wire n_107;
wire n_106;
wire n_105;
wire n_104;
wire n_103;
wire n_102;
wire n_101;
wire n_100;
wire n_99;
wire n_98;
wire n_97;
wire n_96;
wire n_95;
wire n_94;
wire uc_2;


AND2_X1 i_1_125 (.ZN (\Q[31] ), .A1 (n_124), .A2 (i_in2[31]));
MUX2_X1 i_1_124 (.Z (\Q[30] ), .A (i_in2[30]), .B (n_123), .S (i_in2[31]));
MUX2_X1 i_1_123 (.Z (\Q[29] ), .A (i_in2[29]), .B (n_122), .S (i_in2[31]));
MUX2_X1 i_1_122 (.Z (\Q[28] ), .A (i_in2[28]), .B (n_121), .S (i_in2[31]));
MUX2_X1 i_1_121 (.Z (\Q[27] ), .A (i_in2[27]), .B (n_120), .S (i_in2[31]));
MUX2_X1 i_1_120 (.Z (\Q[26] ), .A (i_in2[26]), .B (n_119), .S (i_in2[31]));
MUX2_X1 i_1_119 (.Z (\Q[25] ), .A (i_in2[25]), .B (n_118), .S (i_in2[31]));
MUX2_X1 i_1_118 (.Z (\Q[24] ), .A (i_in2[24]), .B (n_117), .S (i_in2[31]));
MUX2_X1 i_1_117 (.Z (\Q[23] ), .A (i_in2[23]), .B (n_116), .S (i_in2[31]));
MUX2_X1 i_1_116 (.Z (\Q[22] ), .A (i_in2[22]), .B (n_115), .S (i_in2[31]));
MUX2_X1 i_1_115 (.Z (\Q[21] ), .A (i_in2[21]), .B (n_114), .S (i_in2[31]));
MUX2_X1 i_1_114 (.Z (\Q[20] ), .A (i_in2[20]), .B (n_113), .S (i_in2[31]));
MUX2_X1 i_1_113 (.Z (\Q[19] ), .A (i_in2[19]), .B (n_112), .S (i_in2[31]));
MUX2_X1 i_1_112 (.Z (\Q[18] ), .A (i_in2[18]), .B (n_111), .S (i_in2[31]));
MUX2_X1 i_1_111 (.Z (\Q[17] ), .A (i_in2[17]), .B (n_110), .S (i_in2[31]));
MUX2_X1 i_1_110 (.Z (\Q[16] ), .A (i_in2[16]), .B (n_109), .S (i_in2[31]));
MUX2_X1 i_1_109 (.Z (\Q[15] ), .A (i_in2[15]), .B (n_108), .S (i_in2[31]));
MUX2_X1 i_1_108 (.Z (\Q[14] ), .A (i_in2[14]), .B (n_107), .S (i_in2[31]));
MUX2_X1 i_1_107 (.Z (\Q[13] ), .A (i_in2[13]), .B (n_106), .S (i_in2[31]));
MUX2_X1 i_1_106 (.Z (\Q[12] ), .A (i_in2[12]), .B (n_105), .S (i_in2[31]));
MUX2_X1 i_1_105 (.Z (\Q[11] ), .A (i_in2[11]), .B (n_104), .S (i_in2[31]));
MUX2_X1 i_1_104 (.Z (\Q[10] ), .A (i_in2[10]), .B (n_103), .S (i_in2[31]));
MUX2_X1 i_1_103 (.Z (\Q[9] ), .A (i_in2[9]), .B (n_102), .S (i_in2[31]));
MUX2_X1 i_1_102 (.Z (\Q[8] ), .A (i_in2[8]), .B (n_101), .S (i_in2[31]));
MUX2_X1 i_1_101 (.Z (\Q[7] ), .A (i_in2[7]), .B (n_100), .S (i_in2[31]));
MUX2_X1 i_1_100 (.Z (\Q[6] ), .A (i_in2[6]), .B (n_99), .S (i_in2[31]));
MUX2_X1 i_1_99 (.Z (\Q[5] ), .A (i_in2[5]), .B (n_98), .S (i_in2[31]));
MUX2_X1 i_1_98 (.Z (\Q[4] ), .A (i_in2[4]), .B (n_97), .S (i_in2[31]));
MUX2_X1 i_1_97 (.Z (\Q[3] ), .A (i_in2[3]), .B (n_96), .S (i_in2[31]));
MUX2_X1 i_1_96 (.Z (\Q[2] ), .A (i_in2[2]), .B (n_95), .S (i_in2[31]));
MUX2_X1 i_1_95 (.Z (\Q[1] ), .A (i_in2[1]), .B (n_94), .S (i_in2[31]));
AND2_X1 i_1_94 (.ZN (\M[31] ), .A1 (n_93), .A2 (i_in1[31]));
MUX2_X1 i_1_93 (.Z (\M[30] ), .A (i_in1[30]), .B (n_92), .S (i_in1[31]));
MUX2_X1 i_1_92 (.Z (\M[29] ), .A (i_in1[29]), .B (n_91), .S (i_in1[31]));
MUX2_X1 i_1_91 (.Z (\M[28] ), .A (i_in1[28]), .B (n_90), .S (i_in1[31]));
MUX2_X1 i_1_90 (.Z (\M[27] ), .A (i_in1[27]), .B (n_89), .S (i_in1[31]));
MUX2_X1 i_1_89 (.Z (\M[26] ), .A (i_in1[26]), .B (n_88), .S (i_in1[31]));
MUX2_X1 i_1_88 (.Z (\M[25] ), .A (i_in1[25]), .B (n_87), .S (i_in1[31]));
MUX2_X1 i_1_87 (.Z (\M[24] ), .A (i_in1[24]), .B (n_86), .S (i_in1[31]));
MUX2_X1 i_1_86 (.Z (\M[23] ), .A (i_in1[23]), .B (n_85), .S (i_in1[31]));
MUX2_X1 i_1_85 (.Z (\M[22] ), .A (i_in1[22]), .B (n_84), .S (i_in1[31]));
MUX2_X1 i_1_84 (.Z (\M[21] ), .A (i_in1[21]), .B (n_83), .S (i_in1[31]));
MUX2_X1 i_1_83 (.Z (\M[20] ), .A (i_in1[20]), .B (n_82), .S (i_in1[31]));
MUX2_X1 i_1_82 (.Z (\M[19] ), .A (i_in1[19]), .B (n_81), .S (i_in1[31]));
MUX2_X1 i_1_81 (.Z (\M[18] ), .A (i_in1[18]), .B (n_80), .S (i_in1[31]));
MUX2_X1 i_1_80 (.Z (\M[17] ), .A (i_in1[17]), .B (n_79), .S (i_in1[31]));
MUX2_X1 i_1_79 (.Z (\M[16] ), .A (i_in1[16]), .B (n_78), .S (i_in1[31]));
MUX2_X1 i_1_78 (.Z (\M[15] ), .A (i_in1[15]), .B (n_77), .S (i_in1[31]));
MUX2_X1 i_1_77 (.Z (\M[14] ), .A (i_in1[14]), .B (n_76), .S (i_in1[31]));
MUX2_X1 i_1_76 (.Z (\M[13] ), .A (i_in1[13]), .B (n_75), .S (i_in1[31]));
MUX2_X1 i_1_75 (.Z (\M[12] ), .A (i_in1[12]), .B (n_74), .S (i_in1[31]));
MUX2_X1 i_1_74 (.Z (\M[11] ), .A (i_in1[11]), .B (n_73), .S (i_in1[31]));
MUX2_X1 i_1_73 (.Z (\M[10] ), .A (i_in1[10]), .B (n_72), .S (i_in1[31]));
MUX2_X1 i_1_72 (.Z (\M[9] ), .A (i_in1[9]), .B (n_71), .S (i_in1[31]));
MUX2_X1 i_1_71 (.Z (\M[8] ), .A (i_in1[8]), .B (n_70), .S (i_in1[31]));
MUX2_X1 i_1_70 (.Z (\M[7] ), .A (i_in1[7]), .B (n_69), .S (i_in1[31]));
MUX2_X1 i_1_69 (.Z (\M[6] ), .A (i_in1[6]), .B (n_68), .S (i_in1[31]));
MUX2_X1 i_1_68 (.Z (\M[5] ), .A (i_in1[5]), .B (n_67), .S (i_in1[31]));
MUX2_X1 i_1_67 (.Z (\M[4] ), .A (i_in1[4]), .B (n_66), .S (i_in1[31]));
MUX2_X1 i_1_66 (.Z (\M[3] ), .A (i_in1[3]), .B (n_65), .S (i_in1[31]));
MUX2_X1 i_1_65 (.Z (\M[2] ), .A (i_in1[2]), .B (n_64), .S (i_in1[31]));
MUX2_X1 i_1_64 (.Z (\M[1] ), .A (i_in1[1]), .B (n_63), .S (i_in1[31]));
MUX2_X1 i_1_63 (.Z (o_out1[63]), .A (n_62), .B (\out[63] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_62 (.Z (o_out1[62]), .A (n_61), .B (\out[62] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_61 (.Z (o_out1[61]), .A (n_60), .B (\out[61] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_60 (.Z (o_out1[60]), .A (n_59), .B (\out[60] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_59 (.Z (o_out1[59]), .A (n_58), .B (\out[59] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_58 (.Z (o_out1[58]), .A (n_57), .B (\out[58] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_57 (.Z (o_out1[57]), .A (n_56), .B (\out[57] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_56 (.Z (o_out1[56]), .A (n_55), .B (\out[56] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_55 (.Z (o_out1[55]), .A (n_54), .B (\out[55] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_54 (.Z (o_out1[54]), .A (n_53), .B (\out[54] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_53 (.Z (o_out1[53]), .A (n_52), .B (\out[53] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_52 (.Z (o_out1[52]), .A (n_51), .B (\out[52] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_51 (.Z (o_out1[51]), .A (n_50), .B (\out[51] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_50 (.Z (o_out1[50]), .A (n_49), .B (\out[50] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_49 (.Z (o_out1[49]), .A (n_48), .B (\out[49] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_48 (.Z (o_out1[48]), .A (n_47), .B (\out[48] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_47 (.Z (o_out1[47]), .A (n_46), .B (\out[47] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_46 (.Z (o_out1[46]), .A (n_45), .B (\out[46] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_45 (.Z (o_out1[45]), .A (n_44), .B (\out[45] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_44 (.Z (o_out1[44]), .A (n_43), .B (\out[44] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_43 (.Z (o_out1[43]), .A (n_42), .B (\out[43] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_42 (.Z (o_out1[42]), .A (n_41), .B (\out[42] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_41 (.Z (o_out1[41]), .A (n_40), .B (\out[41] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_40 (.Z (o_out1[40]), .A (n_39), .B (\out[40] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_39 (.Z (o_out1[39]), .A (n_38), .B (\out[39] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_38 (.Z (o_out1[38]), .A (n_37), .B (\out[38] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_37 (.Z (o_out1[37]), .A (n_36), .B (\out[37] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_36 (.Z (o_out1[36]), .A (n_35), .B (\out[36] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_35 (.Z (o_out1[35]), .A (n_34), .B (\out[35] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_34 (.Z (o_out1[34]), .A (n_33), .B (\out[34] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_33 (.Z (o_out1[33]), .A (n_32), .B (\out[33] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_32 (.Z (o_out1[32]), .A (n_31), .B (\out[32] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_31 (.Z (o_out1[31]), .A (n_30), .B (\out[31] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_30 (.Z (o_out1[30]), .A (n_29), .B (\out[30] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_29 (.Z (o_out1[29]), .A (n_28), .B (\out[29] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_28 (.Z (o_out1[28]), .A (n_27), .B (\out[28] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_27 (.Z (o_out1[27]), .A (n_26), .B (\out[27] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_26 (.Z (o_out1[26]), .A (n_25), .B (\out[26] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_25 (.Z (o_out1[25]), .A (n_24), .B (\out[25] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_24 (.Z (o_out1[24]), .A (n_23), .B (\out[24] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_23 (.Z (o_out1[23]), .A (n_22), .B (\out[23] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_22 (.Z (o_out1[22]), .A (n_21), .B (\out[22] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_21 (.Z (o_out1[21]), .A (n_20), .B (\out[21] ), .S (hfn_ipo_n5));
MUX2_X1 i_1_20 (.Z (o_out1[20]), .A (n_19), .B (\out[20] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_19 (.Z (o_out1[19]), .A (n_18), .B (\out[19] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_18 (.Z (o_out1[18]), .A (n_17), .B (\out[18] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_17 (.Z (o_out1[17]), .A (n_16), .B (\out[17] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_16 (.Z (o_out1[16]), .A (n_15), .B (\out[16] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_15 (.Z (o_out1[15]), .A (n_14), .B (\out[15] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_14 (.Z (o_out1[14]), .A (n_13), .B (\out[14] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_13 (.Z (o_out1[13]), .A (n_12), .B (\out[13] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_12 (.Z (o_out1[12]), .A (n_11), .B (\out[12] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_11 (.Z (o_out1[11]), .A (n_10), .B (\out[11] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_10 (.Z (o_out1[10]), .A (n_9), .B (\out[10] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_9 (.Z (o_out1[9]), .A (n_8), .B (\out[9] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_8 (.Z (o_out1[8]), .A (n_7), .B (\out[8] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_7 (.Z (o_out1[7]), .A (n_6), .B (\out[7] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_6 (.Z (o_out1[6]), .A (n_5), .B (\out[6] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_5 (.Z (o_out1[5]), .A (n_4), .B (\out[5] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_4 (.Z (o_out1[4]), .A (n_3), .B (\out[4] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_3 (.Z (o_out1[3]), .A (n_2), .B (\out[3] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_2 (.Z (o_out1[2]), .A (n_1), .B (\out[2] ), .S (hfn_ipo_n6));
MUX2_X1 i_1_1 (.Z (o_out1[1]), .A (n_0), .B (\out[1] ), .S (hfn_ipo_n5));
XNOR2_X1 i_1_0 (.ZN (n_1_0), .A (i_in1[31]), .B (i_in2[31]));
datapath__0_26 i_5 (.p_0 ({n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, 
    n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, 
    n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, 
    uc_2}), .i_in2 ({i_in2[31], i_in2[30], i_in2[29], i_in2[28], i_in2[27], i_in2[26], 
    i_in2[25], i_in2[24], i_in2[23], i_in2[22], i_in2[21], i_in2[20], i_in2[19], 
    i_in2[18], i_in2[17], i_in2[16], i_in2[15], i_in2[14], i_in2[13], i_in2[12], 
    i_in2[11], i_in2[10], i_in2[9], i_in2[8], i_in2[7], i_in2[6], i_in2[5], i_in2[4], 
    i_in2[3], i_in2[2], i_in2[1], i_in2[0]}));
datapath__0_24 i_3 (.p_0 ({n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, 
    n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, n_74, n_73, n_72, 
    n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, uc_1}), .i_in1 ({i_in1[31], 
    i_in1[30], i_in1[29], i_in1[28], i_in1[27], i_in1[26], i_in1[25], i_in1[24], 
    i_in1[23], i_in1[22], i_in1[21], i_in1[20], i_in1[19], i_in1[18], i_in1[17], 
    i_in1[16], i_in1[15], i_in1[14], i_in1[13], i_in1[12], i_in1[11], i_in1[10], 
    i_in1[9], i_in1[8], i_in1[7], i_in1[6], i_in1[5], i_in1[4], i_in1[3], i_in1[2], 
    i_in1[1], i_in1[0]}));
datapath__0_21 i_0 (.p_0 ({n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
    n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
    n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, 
    n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, 
    n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, 
    uc_0}), .out ({\out[63] , \out[62] , \out[61] , \out[60] , \out[59] , \out[58] , 
    \out[57] , \out[56] , \out[55] , \out[54] , \out[53] , \out[52] , \out[51] , 
    \out[50] , \out[49] , \out[48] , \out[47] , \out[46] , \out[45] , \out[44] , 
    \out[43] , \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , \out[37] , 
    \out[36] , \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , \out[30] , 
    \out[29] , \out[28] , \out[27] , \out[26] , \out[25] , \out[24] , \out[23] , 
    \out[22] , \out[21] , \out[20] , \out[19] , \out[18] , \out[17] , \out[16] , 
    \out[15] , \out[14] , \out[13] , \out[12] , \out[11] , \out[10] , \out[9] , \out[8] , 
    \out[7] , \out[6] , \out[5] , \out[4] , \out[3] , \out[2] , \out[1] , o_out1[0]}));
shifter shifter (.A ({\A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , 
    \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , 
    \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , 
    \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] }), .o_lsb (lsb), .o_out ({
    \out[63] , \out[62] , \out[61] , \out[60] , \out[59] , \out[58] , \out[57] , 
    \out[56] , \out[55] , \out[54] , \out[53] , \out[52] , \out[51] , \out[50] , 
    \out[49] , \out[48] , \out[47] , \out[46] , \out[45] , \out[44] , \out[43] , 
    \out[42] , \out[41] , \out[40] , \out[39] , \out[38] , \out[37] , \out[36] , 
    \out[35] , \out[34] , \out[33] , \out[32] , \out[31] , \out[30] , \out[29] , 
    \out[28] , \out[27] , \out[26] , \out[25] , \out[24] , \out[23] , \out[22] , 
    \out[21] , \out[20] , \out[19] , \out[18] , \out[17] , \out[16] , \out[15] , 
    \out[14] , \out[13] , \out[12] , \out[11] , \out[10] , \out[9] , \out[8] , \out[7] , 
    \out[6] , \out[5] , \out[4] , \out[3] , \out[2] , \out[1] , o_out1[0]}), .Q ({
    \Q[31] , \Q[30] , \Q[29] , \Q[28] , \Q[27] , \Q[26] , \Q[25] , \Q[24] , \Q[23] , 
    \Q[22] , \Q[21] , \Q[20] , \Q[19] , \Q[18] , \Q[17] , \Q[16] , \Q[15] , \Q[14] , 
    \Q[13] , \Q[12] , \Q[11] , \Q[10] , \Q[9] , \Q[8] , \Q[7] , \Q[6] , \Q[5] , \Q[4] , 
    \Q[3] , \Q[2] , \Q[1] , i_in2[0]}), .i_add (add), .i_adder ({\add_out[32] , \add_out[31] , 
    \add_out[30] , \add_out[29] , \add_out[28] , \add_out[27] , \add_out[26] , \add_out[25] , 
    \add_out[24] , \add_out[23] , \add_out[22] , \add_out[21] , \add_out[20] , \add_out[19] , 
    \add_out[18] , \add_out[17] , \add_out[16] , \add_out[15] , \add_out[14] , \add_out[13] , 
    \add_out[12] , \add_out[11] , \add_out[10] , \add_out[9] , \add_out[8] , \add_out[7] , 
    \add_out[6] , \add_out[5] , \add_out[4] , \add_out[3] , \add_out[2] , \add_out[1] , 
    \add_out[0] }), .i_load (load), .i_out (out_ready), .i_rst (i_rst), .i_shift (shift)
    , .i_clk_CTS_1_PP_0 (CTS_n_tid1_9), .i_clk_CTS_1_PP_1 (i_clk_CTS_1_PP_2));
adder adder (.o_out1 ({\add_out[32] , \add_out[31] , \add_out[30] , \add_out[29] , 
    \add_out[28] , \add_out[27] , \add_out[26] , \add_out[25] , \add_out[24] , \add_out[23] , 
    \add_out[22] , \add_out[21] , \add_out[20] , \add_out[19] , \add_out[18] , \add_out[17] , 
    \add_out[16] , \add_out[15] , \add_out[14] , \add_out[13] , \add_out[12] , \add_out[11] , 
    \add_out[10] , \add_out[9] , \add_out[8] , \add_out[7] , \add_out[6] , \add_out[5] , 
    \add_out[4] , \add_out[3] , \add_out[2] , \add_out[1] , \add_out[0] }), .i_in1 ({
    \M[31] , \M[30] , \M[29] , \M[28] , \M[27] , \M[26] , \M[25] , \M[24] , \M[23] , 
    \M[22] , \M[21] , \M[20] , \M[19] , \M[18] , \M[17] , \M[16] , \M[15] , \M[14] , 
    \M[13] , \M[12] , \M[11] , \M[10] , \M[9] , \M[8] , \M[7] , \M[6] , \M[5] , \M[4] , 
    \M[3] , \M[2] , \M[1] , i_in1[0]}), .i_in2 ({\A[31] , \A[30] , \A[29] , \A[28] , 
    \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , 
    \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , 
    \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] }));
controller controller (.o_add (add), .o_load (load), .o_out (out_ready), .o_shift (shift)
    , .i_clk_CTS_1_PP_0 (CTS_n_tid1_9), .i_lsb (lsb), .i_rst (i_rst), .i_clk_CTS_1_PP_1 (i_clk_CTS_1_PP_0));
CLKBUF_X2 hfn_ipo_c5 (.Z (hfn_ipo_n5), .A (n_1_0));
CLKBUF_X2 hfn_ipo_c6 (.Z (hfn_ipo_n6), .A (n_1_0));

endmodule //multunit

module registerNbits (clk_CTS_1_PP_0, clk_CTS_1_PP_2, clk, reset, en, inp, out);

output [31:0] out;
output clk_CTS_1_PP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_2;
wire drc_ipo_n6;
wire n_0_0;
wire n_1;
wire CTS_n_tid1_8;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CTS_n_tid1_9;
wire CLOCK_slh__n109;
wire CLOCK_slh__n111;
wire CLOCK_slh__n113;
wire CLOCK_slh__n115;
wire CLOCK_slh__n117;
wire CLOCK_slh__n119;
wire CLOCK_slh__n121;
wire CLOCK_slh__n123;
wire CLOCK_slh__n125;
wire CLOCK_slh__n127;
wire CLOCK_slh__n129;
wire CLOCK_slh__n131;
wire CLOCK_slh__n133;
wire CLOCK_slh__n135;
wire CLOCK_slh__n137;
wire CLOCK_slh__n139;
wire CLOCK_slh__n141;
wire CLOCK_slh__n143;
wire CLOCK_slh__n145;
wire CLOCK_slh__n147;
wire CLOCK_slh__n149;
wire CLOCK_slh__n151;
wire CLOCK_slh__n153;
wire CLOCK_slh__n155;
wire CLOCK_slh__n157;
wire CLOCK_slh__n159;
wire CLOCK_slh__n161;
wire CLOCK_slh__n163;
wire CLOCK_slh__n165;
wire CLOCK_slh__n167;
wire CLOCK_slh__n169;
wire CLOCK_slh__n171;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n137), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n169), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n145), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n151), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n139), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n141), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n135), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n131), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n127), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n149), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n117), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n125), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n115), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n147), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n153), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n133), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n129), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n143), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n113), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n123), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n109), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n165), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n111), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n121), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n119), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n163), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n157), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n161), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n167), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n171), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n155), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n159), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (CTS_n_tid1_8), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (CTS_n_tid1_8), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (CTS_n_tid1_8), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (CTS_n_tid1_8), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (CTS_n_tid1_8), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (CTS_n_tid1_8), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (CTS_n_tid1_8), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (CTS_n_tid1_8), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (CTS_n_tid1_8), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (CTS_n_tid1_8), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (CTS_n_tid1_8), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (CTS_n_tid1_8), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (CTS_n_tid1_8), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (CTS_n_tid1_8), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (CTS_n_tid1_8), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (CTS_n_tid1_8), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (CTS_n_tid1_8), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (CTS_n_tid1_8), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (CTS_n_tid1_8), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (CTS_n_tid1_8), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (CTS_n_tid1_8), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (CTS_n_tid1_8), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (CTS_n_tid1_8), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (CTS_n_tid1_8), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (CTS_n_tid1_8), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (CTS_n_tid1_8), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (CTS_n_tid1_8), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (CTS_n_tid1_8), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (CTS_n_tid1_8), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (CTS_n_tid1_8), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (CTS_n_tid1_8), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (CTS_n_tid1_8), .D (n_33));
CLKGATE_X8 clk_gate_out_reg (.GCK (CTS_n_tid1_9), .CK (clk_CTS_1_PP_0), .E (n_1));
BUF_X4 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X3 CTS_L4_c_tid1_6 (.Z (CTS_n_tid1_8), .A (CTS_n_tid1_9));
CLKBUF_X1 CTS_L2_c_tid1_35 (.Z (clk_CTS_1_PP_0), .A (clk_CTS_1_PP_2));
CLKBUF_X1 CLOCK_slh__c42 (.Z (n_13), .A (CLOCK_slh__n109));
CLKBUF_X1 CLOCK_slh__c44 (.Z (n_11), .A (CLOCK_slh__n111));
CLKBUF_X1 CLOCK_slh__c46 (.Z (n_15), .A (CLOCK_slh__n113));
CLKBUF_X1 CLOCK_slh__c48 (.Z (n_21), .A (CLOCK_slh__n115));
CLKBUF_X1 CLOCK_slh__c50 (.Z (n_23), .A (CLOCK_slh__n117));
CLKBUF_X1 CLOCK_slh__c52 (.Z (n_9), .A (CLOCK_slh__n119));
CLKBUF_X1 CLOCK_slh__c54 (.Z (n_10), .A (CLOCK_slh__n121));
CLKBUF_X1 CLOCK_slh__c56 (.Z (n_14), .A (CLOCK_slh__n123));
CLKBUF_X1 CLOCK_slh__c58 (.Z (n_22), .A (CLOCK_slh__n125));
CLKBUF_X1 CLOCK_slh__c60 (.Z (n_25), .A (CLOCK_slh__n127));
CLKBUF_X1 CLOCK_slh__c62 (.Z (n_17), .A (CLOCK_slh__n129));
CLKBUF_X1 CLOCK_slh__c64 (.Z (n_26), .A (CLOCK_slh__n131));
CLKBUF_X1 CLOCK_slh__c66 (.Z (n_18), .A (CLOCK_slh__n133));
CLKBUF_X1 CLOCK_slh__c68 (.Z (n_27), .A (CLOCK_slh__n135));
CLKBUF_X1 CLOCK_slh__c70 (.Z (n_33), .A (CLOCK_slh__n137));
CLKBUF_X1 CLOCK_slh__c72 (.Z (n_29), .A (CLOCK_slh__n139));
CLKBUF_X1 CLOCK_slh__c74 (.Z (n_28), .A (CLOCK_slh__n141));
CLKBUF_X1 CLOCK_slh__c76 (.Z (n_16), .A (CLOCK_slh__n143));
CLKBUF_X1 CLOCK_slh__c78 (.Z (n_31), .A (CLOCK_slh__n145));
CLKBUF_X1 CLOCK_slh__c80 (.Z (n_20), .A (CLOCK_slh__n147));
CLKBUF_X1 CLOCK_slh__c82 (.Z (n_24), .A (CLOCK_slh__n149));
CLKBUF_X1 CLOCK_slh__c84 (.Z (n_30), .A (CLOCK_slh__n151));
CLKBUF_X1 CLOCK_slh__c86 (.Z (n_19), .A (CLOCK_slh__n153));
CLKBUF_X1 CLOCK_slh__c88 (.Z (n_3), .A (CLOCK_slh__n155));
CLKBUF_X1 CLOCK_slh__c90 (.Z (n_7), .A (CLOCK_slh__n157));
CLKBUF_X1 CLOCK_slh__c92 (.Z (n_2), .A (CLOCK_slh__n159));
CLKBUF_X1 CLOCK_slh__c94 (.Z (n_6), .A (CLOCK_slh__n161));
CLKBUF_X1 CLOCK_slh__c96 (.Z (n_8), .A (CLOCK_slh__n163));
CLKBUF_X1 CLOCK_slh__c98 (.Z (n_12), .A (CLOCK_slh__n165));
CLKBUF_X1 CLOCK_slh__c100 (.Z (n_5), .A (CLOCK_slh__n167));
CLKBUF_X1 CLOCK_slh__c102 (.Z (n_32), .A (CLOCK_slh__n169));
CLKBUF_X1 CLOCK_slh__c104 (.Z (n_4), .A (CLOCK_slh__n171));

endmodule //registerNbits

module registerNbits__0_32 (clk_CTS_1_PP_0, clk_CTS_1_PP_1, clk, reset, en, inp, 
    out);

output [31:0] out;
output clk_CTS_1_PP_0;
input clk;
input en;
input [31:0] inp;
input reset;
input clk_CTS_1_PP_1;
wire drc_ipo_n6;
wire n_0_0;
wire n_1;
wire n_0;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_25;
wire n_24;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;
wire CLOCK_slh__n65;
wire CLOCK_slh__n67;
wire CLOCK_slh__n69;
wire CLOCK_slh__n71;
wire CLOCK_slh__n73;
wire CLOCK_slh__n75;
wire CLOCK_slh__n77;
wire CLOCK_slh__n79;
wire CLOCK_slh__n81;
wire CLOCK_slh__n83;
wire CLOCK_slh__n85;
wire CLOCK_slh__n87;
wire CLOCK_slh__n89;
wire CLOCK_slh__n91;
wire CLOCK_slh__n93;
wire CLOCK_slh__n95;
wire CLOCK_slh__n97;
wire CLOCK_slh__n99;
wire CLOCK_slh__n101;
wire CLOCK_slh__n103;
wire CLOCK_slh__n105;
wire CLOCK_slh__n107;
wire CLOCK_slh__n108;
wire CLOCK_slh__n109;
wire CLOCK_slh__n110;
wire CLOCK_slh__n111;
wire CLOCK_slh__n112;
wire CLOCK_slh__n113;
wire CLOCK_slh__n114;
wire CLOCK_slh__n115;
wire CLOCK_slh__n116;
wire CLOCK_slh__n117;


AND2_X1 i_0_33 (.ZN (CLOCK_slh__n71), .A1 (n_0_0), .A2 (inp[31]));
AND2_X1 i_0_32 (.ZN (CLOCK_slh__n69), .A1 (n_0_0), .A2 (inp[30]));
AND2_X1 i_0_31 (.ZN (CLOCK_slh__n73), .A1 (n_0_0), .A2 (inp[29]));
AND2_X1 i_0_30 (.ZN (CLOCK_slh__n93), .A1 (n_0_0), .A2 (inp[28]));
AND2_X1 i_0_29 (.ZN (CLOCK_slh__n75), .A1 (n_0_0), .A2 (inp[27]));
AND2_X1 i_0_28 (.ZN (CLOCK_slh__n65), .A1 (n_0_0), .A2 (inp[26]));
AND2_X1 i_0_27 (.ZN (CLOCK_slh__n91), .A1 (n_0_0), .A2 (inp[25]));
AND2_X1 i_0_26 (.ZN (CLOCK_slh__n101), .A1 (n_0_0), .A2 (inp[24]));
AND2_X1 i_0_25 (.ZN (CLOCK_slh__n83), .A1 (n_0_0), .A2 (inp[23]));
AND2_X1 i_0_24 (.ZN (CLOCK_slh__n99), .A1 (n_0_0), .A2 (inp[22]));
AND2_X1 i_0_23 (.ZN (CLOCK_slh__n81), .A1 (n_0_0), .A2 (inp[21]));
AND2_X1 i_0_22 (.ZN (CLOCK_slh__n77), .A1 (n_0_0), .A2 (inp[20]));
AND2_X1 i_0_21 (.ZN (CLOCK_slh__n95), .A1 (n_0_0), .A2 (inp[19]));
AND2_X1 i_0_20 (.ZN (CLOCK_slh__n97), .A1 (n_0_0), .A2 (inp[18]));
AND2_X1 i_0_19 (.ZN (CLOCK_slh__n67), .A1 (n_0_0), .A2 (inp[17]));
AND2_X1 i_0_18 (.ZN (CLOCK_slh__n107), .A1 (n_0_0), .A2 (inp[16]));
AND2_X1 i_0_17 (.ZN (CLOCK_slh__n79), .A1 (n_0_0), .A2 (inp[15]));
AND2_X1 i_0_16 (.ZN (CLOCK_slh__n87), .A1 (n_0_0), .A2 (inp[14]));
AND2_X1 i_0_15 (.ZN (CLOCK_slh__n85), .A1 (n_0_0), .A2 (inp[13]));
AND2_X1 i_0_14 (.ZN (CLOCK_slh__n89), .A1 (n_0_0), .A2 (inp[12]));
AND2_X1 i_0_13 (.ZN (CLOCK_slh__n105), .A1 (n_0_0), .A2 (inp[11]));
AND2_X1 i_0_12 (.ZN (CLOCK_slh__n103), .A1 (n_0_0), .A2 (inp[10]));
AND2_X1 i_0_11 (.ZN (CLOCK_slh__n109), .A1 (n_0_0), .A2 (inp[9]));
AND2_X1 i_0_10 (.ZN (CLOCK_slh__n108), .A1 (n_0_0), .A2 (inp[8]));
AND2_X1 i_0_9 (.ZN (CLOCK_slh__n110), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (CLOCK_slh__n111), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (CLOCK_slh__n113), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (CLOCK_slh__n115), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (CLOCK_slh__n117), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (CLOCK_slh__n116), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (CLOCK_slh__n112), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (CLOCK_slh__n114), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
DFF_X1 \out_reg[8]  (.Q (out[8]), .CK (n_0), .D (n_10));
DFF_X1 \out_reg[9]  (.Q (out[9]), .CK (n_0), .D (n_11));
DFF_X1 \out_reg[10]  (.Q (out[10]), .CK (n_0), .D (n_12));
DFF_X1 \out_reg[11]  (.Q (out[11]), .CK (n_0), .D (n_13));
DFF_X1 \out_reg[12]  (.Q (out[12]), .CK (n_0), .D (n_14));
DFF_X1 \out_reg[13]  (.Q (out[13]), .CK (n_0), .D (n_15));
DFF_X1 \out_reg[14]  (.Q (out[14]), .CK (n_0), .D (n_16));
DFF_X1 \out_reg[15]  (.Q (out[15]), .CK (n_0), .D (n_17));
DFF_X1 \out_reg[16]  (.Q (out[16]), .CK (n_0), .D (n_18));
DFF_X1 \out_reg[17]  (.Q (out[17]), .CK (n_0), .D (n_19));
DFF_X1 \out_reg[18]  (.Q (out[18]), .CK (n_0), .D (n_20));
DFF_X1 \out_reg[19]  (.Q (out[19]), .CK (n_0), .D (n_21));
DFF_X1 \out_reg[20]  (.Q (out[20]), .CK (n_0), .D (n_22));
DFF_X1 \out_reg[21]  (.Q (out[21]), .CK (n_0), .D (n_23));
DFF_X1 \out_reg[22]  (.Q (out[22]), .CK (n_0), .D (n_24));
DFF_X1 \out_reg[23]  (.Q (out[23]), .CK (n_0), .D (n_25));
DFF_X1 \out_reg[24]  (.Q (out[24]), .CK (n_0), .D (n_26));
DFF_X1 \out_reg[25]  (.Q (out[25]), .CK (n_0), .D (n_27));
DFF_X1 \out_reg[26]  (.Q (out[26]), .CK (n_0), .D (n_28));
DFF_X1 \out_reg[27]  (.Q (out[27]), .CK (n_0), .D (n_29));
DFF_X1 \out_reg[28]  (.Q (out[28]), .CK (n_0), .D (n_30));
DFF_X1 \out_reg[29]  (.Q (out[29]), .CK (n_0), .D (n_31));
DFF_X1 \out_reg[30]  (.Q (out[30]), .CK (n_0), .D (n_32));
DFF_X1 \out_reg[31]  (.Q (drc_ipo_n6), .CK (n_0), .D (n_33));
CLKGATE_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk_CTS_1_PP_0), .E (n_1));
BUF_X4 drc_ipo_c3 (.Z (out[31]), .A (drc_ipo_n6));
CLKBUF_X3 CTS_L1_c_tid1_10 (.Z (clk_CTS_1_PP_0), .A (clk_CTS_1_PP_1));
CLKBUF_X1 CLOCK_slh__c17 (.Z (n_28), .A (CLOCK_slh__n65));
CLKBUF_X1 CLOCK_slh__c19 (.Z (n_19), .A (CLOCK_slh__n67));
CLKBUF_X1 CLOCK_slh__c21 (.Z (n_32), .A (CLOCK_slh__n69));
CLKBUF_X1 CLOCK_slh__c23 (.Z (n_33), .A (CLOCK_slh__n71));
CLKBUF_X1 CLOCK_slh__c25 (.Z (n_31), .A (CLOCK_slh__n73));
CLKBUF_X1 CLOCK_slh__c27 (.Z (n_29), .A (CLOCK_slh__n75));
CLKBUF_X1 CLOCK_slh__c29 (.Z (n_22), .A (CLOCK_slh__n77));
CLKBUF_X1 CLOCK_slh__c31 (.Z (n_17), .A (CLOCK_slh__n79));
CLKBUF_X1 CLOCK_slh__c33 (.Z (n_23), .A (CLOCK_slh__n81));
CLKBUF_X1 CLOCK_slh__c35 (.Z (n_25), .A (CLOCK_slh__n83));
CLKBUF_X1 CLOCK_slh__c37 (.Z (n_15), .A (CLOCK_slh__n85));
CLKBUF_X1 CLOCK_slh__c39 (.Z (n_16), .A (CLOCK_slh__n87));
CLKBUF_X1 CLOCK_slh__c41 (.Z (n_14), .A (CLOCK_slh__n89));
CLKBUF_X1 CLOCK_slh__c43 (.Z (n_27), .A (CLOCK_slh__n91));
CLKBUF_X1 CLOCK_slh__c45 (.Z (n_30), .A (CLOCK_slh__n93));
CLKBUF_X1 CLOCK_slh__c47 (.Z (n_21), .A (CLOCK_slh__n95));
CLKBUF_X1 CLOCK_slh__c49 (.Z (n_20), .A (CLOCK_slh__n97));
CLKBUF_X1 CLOCK_slh__c51 (.Z (n_24), .A (CLOCK_slh__n99));
CLKBUF_X1 CLOCK_slh__c53 (.Z (n_26), .A (CLOCK_slh__n101));
CLKBUF_X1 CLOCK_slh__c55 (.Z (n_12), .A (CLOCK_slh__n103));
CLKBUF_X1 CLOCK_slh__c57 (.Z (n_13), .A (CLOCK_slh__n105));
CLKBUF_X1 CLOCK_slh__c59 (.Z (n_18), .A (CLOCK_slh__n107));
CLKBUF_X1 CLOCK_slh__c60 (.Z (n_10), .A (CLOCK_slh__n108));
CLKBUF_X1 CLOCK_slh__c61 (.Z (n_11), .A (CLOCK_slh__n109));
CLKBUF_X1 CLOCK_slh__c62 (.Z (n_9), .A (CLOCK_slh__n110));
CLKBUF_X1 CLOCK_slh__c63 (.Z (n_8), .A (CLOCK_slh__n111));
CLKBUF_X1 CLOCK_slh__c64 (.Z (n_3), .A (CLOCK_slh__n112));
CLKBUF_X1 CLOCK_slh__c65 (.Z (n_7), .A (CLOCK_slh__n113));
CLKBUF_X1 CLOCK_slh__c66 (.Z (n_2), .A (CLOCK_slh__n114));
CLKBUF_X1 CLOCK_slh__c67 (.Z (n_6), .A (CLOCK_slh__n115));
CLKBUF_X1 CLOCK_slh__c68 (.Z (n_4), .A (CLOCK_slh__n116));
CLKBUF_X1 CLOCK_slh__c69 (.Z (n_5), .A (CLOCK_slh__n117));

endmodule //registerNbits__0_32

module sequential (i_clk, i_rst, i_en, i_inputA, i_inputB, o_result);

output [63:0] o_result;
input i_clk;
input i_en;
input [31:0] i_inputA;
input [31:0] i_inputB;
input i_rst;
wire CTS_n_tid1_3;
wire \A_reg[31] ;
wire \A_reg[30] ;
wire \A_reg[29] ;
wire \A_reg[28] ;
wire \A_reg[27] ;
wire \A_reg[26] ;
wire \A_reg[25] ;
wire \A_reg[24] ;
wire \A_reg[23] ;
wire \A_reg[22] ;
wire \A_reg[21] ;
wire \A_reg[20] ;
wire \A_reg[19] ;
wire \A_reg[18] ;
wire \A_reg[17] ;
wire \A_reg[16] ;
wire \A_reg[15] ;
wire \A_reg[14] ;
wire \A_reg[13] ;
wire \A_reg[12] ;
wire \A_reg[11] ;
wire \A_reg[10] ;
wire \A_reg[9] ;
wire \A_reg[8] ;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[31] ;
wire \B_reg[30] ;
wire \B_reg[29] ;
wire \B_reg[28] ;
wire \B_reg[27] ;
wire \B_reg[26] ;
wire \B_reg[25] ;
wire \B_reg[24] ;
wire \B_reg[23] ;
wire \B_reg[22] ;
wire \B_reg[21] ;
wire \B_reg[20] ;
wire \B_reg[19] ;
wire \B_reg[18] ;
wire \B_reg[17] ;
wire \B_reg[16] ;
wire \B_reg[15] ;
wire \B_reg[14] ;
wire \B_reg[13] ;
wire \B_reg[12] ;
wire \B_reg[11] ;
wire \B_reg[10] ;
wire \B_reg[9] ;
wire \B_reg[8] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire \out_reg[63] ;
wire \out_reg[62] ;
wire \out_reg[61] ;
wire \out_reg[60] ;
wire \out_reg[59] ;
wire \out_reg[58] ;
wire \out_reg[57] ;
wire \out_reg[56] ;
wire \out_reg[55] ;
wire \out_reg[54] ;
wire \out_reg[53] ;
wire \out_reg[52] ;
wire \out_reg[51] ;
wire \out_reg[50] ;
wire \out_reg[49] ;
wire \out_reg[48] ;
wire \out_reg[47] ;
wire \out_reg[46] ;
wire \out_reg[45] ;
wire \out_reg[44] ;
wire \out_reg[43] ;
wire \out_reg[42] ;
wire \out_reg[41] ;
wire \out_reg[40] ;
wire \out_reg[39] ;
wire \out_reg[38] ;
wire \out_reg[37] ;
wire \out_reg[36] ;
wire \out_reg[35] ;
wire \out_reg[34] ;
wire \out_reg[33] ;
wire \out_reg[32] ;
wire \out_reg[31] ;
wire \out_reg[30] ;
wire \out_reg[29] ;
wire \out_reg[28] ;
wire \out_reg[27] ;
wire \out_reg[26] ;
wire \out_reg[25] ;
wire \out_reg[24] ;
wire \out_reg[23] ;
wire \out_reg[22] ;
wire \out_reg[21] ;
wire \out_reg[20] ;
wire \out_reg[19] ;
wire \out_reg[18] ;
wire \out_reg[17] ;
wire \out_reg[16] ;
wire \out_reg[15] ;
wire \out_reg[14] ;
wire \out_reg[13] ;
wire \out_reg[12] ;
wire \out_reg[11] ;
wire \out_reg[10] ;
wire \out_reg[9] ;
wire \out_reg[8] ;
wire \out_reg[7] ;
wire \out_reg[6] ;
wire \out_reg[5] ;
wire \out_reg[4] ;
wire \out_reg[3] ;
wire \out_reg[2] ;
wire \out_reg[1] ;
wire \out_reg[0] ;
wire CTS_n_tid1_7;


registerNbits__parameterized0 outReg (.out ({o_result[63], o_result[62], o_result[61], 
    o_result[60], o_result[59], o_result[58], o_result[57], o_result[56], o_result[55], 
    o_result[54], o_result[53], o_result[52], o_result[51], o_result[50], o_result[49], 
    o_result[48], o_result[47], o_result[46], o_result[45], o_result[44], o_result[43], 
    o_result[42], o_result[41], o_result[40], o_result[39], o_result[38], o_result[37], 
    o_result[36], o_result[35], o_result[34], o_result[33], o_result[32], o_result[31], 
    o_result[30], o_result[29], o_result[28], o_result[27], o_result[26], o_result[25], 
    o_result[24], o_result[23], o_result[22], o_result[21], o_result[20], o_result[19], 
    o_result[18], o_result[17], o_result[16], o_result[15], o_result[14], o_result[13], 
    o_result[12], o_result[11], o_result[10], o_result[9], o_result[8], o_result[7], 
    o_result[6], o_result[5], o_result[4], o_result[3], o_result[2], o_result[1], 
    o_result[0]}), .en (i_en), .inp ({\out_reg[63] , \out_reg[62] , \out_reg[61] , 
    \out_reg[60] , \out_reg[59] , \out_reg[58] , \out_reg[57] , \out_reg[56] , \out_reg[55] , 
    \out_reg[54] , \out_reg[53] , \out_reg[52] , \out_reg[51] , \out_reg[50] , \out_reg[49] , 
    \out_reg[48] , \out_reg[47] , \out_reg[46] , \out_reg[45] , \out_reg[44] , \out_reg[43] , 
    \out_reg[42] , \out_reg[41] , \out_reg[40] , \out_reg[39] , \out_reg[38] , \out_reg[37] , 
    \out_reg[36] , \out_reg[35] , \out_reg[34] , \out_reg[33] , \out_reg[32] , \out_reg[31] , 
    \out_reg[30] , \out_reg[29] , \out_reg[28] , \out_reg[27] , \out_reg[26] , \out_reg[25] , 
    \out_reg[24] , \out_reg[23] , \out_reg[22] , \out_reg[21] , \out_reg[20] , \out_reg[19] , 
    \out_reg[18] , \out_reg[17] , \out_reg[16] , \out_reg[15] , \out_reg[14] , \out_reg[13] , 
    \out_reg[12] , \out_reg[11] , \out_reg[10] , \out_reg[9] , \out_reg[8] , \out_reg[7] , 
    \out_reg[6] , \out_reg[5] , \out_reg[4] , \out_reg[3] , \out_reg[2] , \out_reg[1] , 
    \out_reg[0] }), .reset (i_rst), .clk_CTS_1_PP_0 (CTS_n_tid1_7));
multunit mult (.o_out1 ({\out_reg[63] , \out_reg[62] , \out_reg[61] , \out_reg[60] , 
    \out_reg[59] , \out_reg[58] , \out_reg[57] , \out_reg[56] , \out_reg[55] , \out_reg[54] , 
    \out_reg[53] , \out_reg[52] , \out_reg[51] , \out_reg[50] , \out_reg[49] , \out_reg[48] , 
    \out_reg[47] , \out_reg[46] , \out_reg[45] , \out_reg[44] , \out_reg[43] , \out_reg[42] , 
    \out_reg[41] , \out_reg[40] , \out_reg[39] , \out_reg[38] , \out_reg[37] , \out_reg[36] , 
    \out_reg[35] , \out_reg[34] , \out_reg[33] , \out_reg[32] , \out_reg[31] , \out_reg[30] , 
    \out_reg[29] , \out_reg[28] , \out_reg[27] , \out_reg[26] , \out_reg[25] , \out_reg[24] , 
    \out_reg[23] , \out_reg[22] , \out_reg[21] , \out_reg[20] , \out_reg[19] , \out_reg[18] , 
    \out_reg[17] , \out_reg[16] , \out_reg[15] , \out_reg[14] , \out_reg[13] , \out_reg[12] , 
    \out_reg[11] , \out_reg[10] , \out_reg[9] , \out_reg[8] , \out_reg[7] , \out_reg[6] , 
    \out_reg[5] , \out_reg[4] , \out_reg[3] , \out_reg[2] , \out_reg[1] , \out_reg[0] })
    , .i_in1 ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , \A_reg[27] , \A_reg[26] , 
    \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , \A_reg[21] , \A_reg[20] , 
    \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , \A_reg[15] , \A_reg[14] , 
    \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , \A_reg[9] , \A_reg[8] , \A_reg[7] , 
    \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , \A_reg[1] , \A_reg[0] })
    , .i_in2 ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , \B_reg[26] , 
    \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , \B_reg[20] , 
    \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , \B_reg[14] , 
    \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , \B_reg[8] , \B_reg[7] , 
    \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] })
    , .i_rst (i_rst), .i_clk_CTS_1_PP_0 (CTS_n_tid1_3), .i_clk_CTS_1_PP_2 (CTS_n_tid1_7));
registerNbits regB (.out ({\B_reg[31] , \B_reg[30] , \B_reg[29] , \B_reg[28] , \B_reg[27] , 
    \B_reg[26] , \B_reg[25] , \B_reg[24] , \B_reg[23] , \B_reg[22] , \B_reg[21] , 
    \B_reg[20] , \B_reg[19] , \B_reg[18] , \B_reg[17] , \B_reg[16] , \B_reg[15] , 
    \B_reg[14] , \B_reg[13] , \B_reg[12] , \B_reg[11] , \B_reg[10] , \B_reg[9] , 
    \B_reg[8] , \B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , \B_reg[2] , 
    \B_reg[1] , \B_reg[0] }), .clk_CTS_1_PP_0 (CTS_n_tid1_3), .en (i_en), .inp ({
    i_inputB[31], i_inputB[30], i_inputB[29], i_inputB[28], i_inputB[27], i_inputB[26], 
    i_inputB[25], i_inputB[24], i_inputB[23], i_inputB[22], i_inputB[21], i_inputB[20], 
    i_inputB[19], i_inputB[18], i_inputB[17], i_inputB[16], i_inputB[15], i_inputB[14], 
    i_inputB[13], i_inputB[12], i_inputB[11], i_inputB[10], i_inputB[9], i_inputB[8], 
    i_inputB[7], i_inputB[6], i_inputB[5], i_inputB[4], i_inputB[3], i_inputB[2], 
    i_inputB[1], i_inputB[0]}), .reset (i_rst), .clk_CTS_1_PP_2 (CTS_n_tid1_7));
registerNbits__0_32 regA (.out ({\A_reg[31] , \A_reg[30] , \A_reg[29] , \A_reg[28] , 
    \A_reg[27] , \A_reg[26] , \A_reg[25] , \A_reg[24] , \A_reg[23] , \A_reg[22] , 
    \A_reg[21] , \A_reg[20] , \A_reg[19] , \A_reg[18] , \A_reg[17] , \A_reg[16] , 
    \A_reg[15] , \A_reg[14] , \A_reg[13] , \A_reg[12] , \A_reg[11] , \A_reg[10] , 
    \A_reg[9] , \A_reg[8] , \A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .clk_CTS_1_PP_0 (CTS_n_tid1_7), .en (i_en)
    , .inp ({i_inputA[31], i_inputA[30], i_inputA[29], i_inputA[28], i_inputA[27], 
    i_inputA[26], i_inputA[25], i_inputA[24], i_inputA[23], i_inputA[22], i_inputA[21], 
    i_inputA[20], i_inputA[19], i_inputA[18], i_inputA[17], i_inputA[16], i_inputA[15], 
    i_inputA[14], i_inputA[13], i_inputA[12], i_inputA[11], i_inputA[10], i_inputA[9], 
    i_inputA[8], i_inputA[7], i_inputA[6], i_inputA[5], i_inputA[4], i_inputA[3], 
    i_inputA[2], i_inputA[1], i_inputA[0]}), .reset (i_rst), .clk_CTS_1_PP_1 (i_clk));

endmodule //sequential


