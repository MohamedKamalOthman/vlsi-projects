/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Nov  2 22:14:20 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1112292000 */

module halfAdder__0_300(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_301(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_300 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_292(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_289(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_293(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_292 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_289 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_284(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_281(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_285(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_284 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_281 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_276(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_273(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_277(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_276 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_273 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_268(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_265(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_269(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_268 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_265 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_260(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_257(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_261(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_260 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_257 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_252(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_249(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_253(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_252 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_249 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_244(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_241(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_245(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_244 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_241 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_236(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_233(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_237(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_236 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_233 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_228(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_225(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_229(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_228 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_225 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_220(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_217(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_221(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_220 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_217 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_212(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_209(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_213(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_212 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_209 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_204(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_201(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_205(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_204 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_201 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_196(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_193(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_197(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_196 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_193 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_188(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_185(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_189(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_188 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_185 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_180(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_177(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_181(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_180 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_177 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module __RippleAdder____0_302(cin, x, y, cout, sum);
   input cin;
   input [15:0]x;
   input [15:0]y;
   output cout;
   output [15:0]sum;

   wire [14:0]coutWires;

   fullAdder__0_301 genblk1_0_FA (.cin(), .x(x[0]), .y(y[0]), .cout(coutWires[0]), 
      .sum(sum[0]));
   fullAdder__0_293 genblk1_1_FA3 (.cin(coutWires[0]), .x(x[1]), .y(y[1]), 
      .cout(coutWires[1]), .sum(sum[1]));
   fullAdder__0_285 genblk1_2_FA3 (.cin(coutWires[1]), .x(x[2]), .y(y[2]), 
      .cout(coutWires[2]), .sum(sum[2]));
   fullAdder__0_277 genblk1_3_FA3 (.cin(coutWires[2]), .x(x[3]), .y(y[3]), 
      .cout(coutWires[3]), .sum(sum[3]));
   fullAdder__0_269 genblk1_4_FA3 (.cin(coutWires[3]), .x(x[4]), .y(y[4]), 
      .cout(coutWires[4]), .sum(sum[4]));
   fullAdder__0_261 genblk1_5_FA3 (.cin(coutWires[4]), .x(x[5]), .y(y[5]), 
      .cout(coutWires[5]), .sum(sum[5]));
   fullAdder__0_253 genblk1_6_FA3 (.cin(coutWires[5]), .x(x[6]), .y(y[6]), 
      .cout(coutWires[6]), .sum(sum[6]));
   fullAdder__0_245 genblk1_7_FA3 (.cin(coutWires[6]), .x(x[7]), .y(y[7]), 
      .cout(coutWires[7]), .sum(sum[7]));
   fullAdder__0_237 genblk1_8_FA3 (.cin(coutWires[7]), .x(x[8]), .y(y[8]), 
      .cout(coutWires[8]), .sum(sum[8]));
   fullAdder__0_229 genblk1_9_FA3 (.cin(coutWires[8]), .x(x[9]), .y(y[9]), 
      .cout(coutWires[9]), .sum(sum[9]));
   fullAdder__0_221 genblk1_10_FA3 (.cin(coutWires[9]), .x(x[10]), .y(y[10]), 
      .cout(coutWires[10]), .sum(sum[10]));
   fullAdder__0_213 genblk1_11_FA3 (.cin(coutWires[10]), .x(x[11]), .y(y[11]), 
      .cout(coutWires[11]), .sum(sum[11]));
   fullAdder__0_205 genblk1_12_FA3 (.cin(coutWires[11]), .x(x[12]), .y(y[12]), 
      .cout(coutWires[12]), .sum(sum[12]));
   fullAdder__0_197 genblk1_13_FA3 (.cin(coutWires[12]), .x(x[13]), .y(y[13]), 
      .cout(coutWires[13]), .sum(sum[13]));
   fullAdder__0_189 genblk1_14_FA3 (.cin(coutWires[13]), .x(x[14]), .y(y[14]), 
      .cout(coutWires[14]), .sum(sum[14]));
   fullAdder__0_181 genblk1_15_FA2 (.cin(coutWires[14]), .x(x[15]), .y(y[15]), 
      .cout(cout), .sum(sum[15]));
endmodule

module halfAdder__0_60(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_61(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_60 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_68(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_65(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_69(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_68 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_65 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_76(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_73(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_77(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_76 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_73 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_84(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_81(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_85(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_84 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_81 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_92(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_89(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_93(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_92 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_89 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_100(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_97(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_101(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_100 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_97 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_108(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_105(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_109(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_108 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_105 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_116(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_113(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_117(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_116 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_113 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_124(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_121(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_125(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_124 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_121 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_132(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_129(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_133(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_132 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_129 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_140(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_137(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_141(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_140 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_137 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_148(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_145(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_149(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_148 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_145 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_156(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_153(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_157(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_156 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_153 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_164(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_161(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_165(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_164 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_161 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_172(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_169(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_173(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_172 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_169 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_5(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_8(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_5 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_8 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module __RippleAdder__(cin, x, y, cout, sum);
   input cin;
   input [15:0]x;
   input [15:0]y;
   output cout;
   output [15:0]sum;

   wire [14:0]coutWires;

   fullAdder__0_61 genblk1_0_FA (.cin(), .x(x[0]), .y(y[0]), .cout(coutWires[0]), 
      .sum(sum[0]));
   fullAdder__0_69 genblk1_1_FA3 (.cin(coutWires[0]), .x(x[1]), .y(y[1]), 
      .cout(coutWires[1]), .sum(sum[1]));
   fullAdder__0_77 genblk1_2_FA3 (.cin(coutWires[1]), .x(x[2]), .y(y[2]), 
      .cout(coutWires[2]), .sum(sum[2]));
   fullAdder__0_85 genblk1_3_FA3 (.cin(coutWires[2]), .x(x[3]), .y(y[3]), 
      .cout(coutWires[3]), .sum(sum[3]));
   fullAdder__0_93 genblk1_4_FA3 (.cin(coutWires[3]), .x(x[4]), .y(y[4]), 
      .cout(coutWires[4]), .sum(sum[4]));
   fullAdder__0_101 genblk1_5_FA3 (.cin(coutWires[4]), .x(x[5]), .y(y[5]), 
      .cout(coutWires[5]), .sum(sum[5]));
   fullAdder__0_109 genblk1_6_FA3 (.cin(coutWires[5]), .x(x[6]), .y(y[6]), 
      .cout(coutWires[6]), .sum(sum[6]));
   fullAdder__0_117 genblk1_7_FA3 (.cin(coutWires[6]), .x(x[7]), .y(y[7]), 
      .cout(coutWires[7]), .sum(sum[7]));
   fullAdder__0_125 genblk1_8_FA3 (.cin(coutWires[7]), .x(x[8]), .y(y[8]), 
      .cout(coutWires[8]), .sum(sum[8]));
   fullAdder__0_133 genblk1_9_FA3 (.cin(coutWires[8]), .x(x[9]), .y(y[9]), 
      .cout(coutWires[9]), .sum(sum[9]));
   fullAdder__0_141 genblk1_10_FA3 (.cin(coutWires[9]), .x(x[10]), .y(y[10]), 
      .cout(coutWires[10]), .sum(sum[10]));
   fullAdder__0_149 genblk1_11_FA3 (.cin(coutWires[10]), .x(x[11]), .y(y[11]), 
      .cout(coutWires[11]), .sum(sum[11]));
   fullAdder__0_157 genblk1_12_FA3 (.cin(coutWires[11]), .x(x[12]), .y(y[12]), 
      .cout(coutWires[12]), .sum(sum[12]));
   fullAdder__0_165 genblk1_13_FA3 (.cin(coutWires[12]), .x(x[13]), .y(y[13]), 
      .cout(coutWires[13]), .sum(sum[13]));
   fullAdder__0_173 genblk1_14_FA3 (.cin(coutWires[13]), .x(x[14]), .y(y[14]), 
      .cout(coutWires[14]), .sum(sum[14]));
   fullAdder genblk1_15_FA2 (.cin(coutWires[14]), .x(x[15]), .y(y[15]), .cout(
      cout), .sum(sum[15]));
endmodule

module halfAdder__0_11(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_14(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_17(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_20(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_23(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_26(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_29(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_32(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_35(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_38(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_41(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_44(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_47(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_50(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_53(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module carryIncrementAdder(in1, in2, sum);
   input [31:0]in1;
   input [31:0]in2;
   output [32:0]sum;

   wire coutWire;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire carryWires;

   __RippleAdder____0_302 RA1 (.cin(), .x({in1[15], in1[14], in1[13], in1[12], 
      in1[11], in1[10], in1[9], in1[8], in1[7], in1[6], in1[5], in1[4], in1[3], 
      in1[2], in1[1], in1[0]}), .y({in2[15], in2[14], in2[13], in2[12], in2[11], 
      in2[10], in2[9], in2[8], in2[7], in2[6], in2[5], in2[4], in2[3], in2[2], 
      in2[1], in2[0]}), .cout(coutWire), .sum({sum[15], sum[14], sum[13], 
      sum[12], sum[11], sum[10], sum[9], sum[8], sum[7], sum[6], sum[5], sum[4], 
      sum[3], sum[2], sum[1], sum[0]}));
   __RippleAdder__ RA2 (.cin(), .x({in1[31], in1[30], in1[29], in1[28], in1[27], 
      in1[26], in1[25], in1[24], in1[23], in1[22], in1[21], in1[20], in1[19], 
      in1[18], in1[17], in1[16]}), .y({in2[31], in2[30], in2[29], in2[28], 
      in2[27], in2[26], in2[25], in2[24], in2[23], in2[22], in2[21], in2[20], 
      in2[19], in2[18], in2[17], in2[16]}), .cout(n_0_16), .sum({n_0_15, n_0_14, 
      n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
      n_0_3, n_0_2, n_0_1, n_0_0}));
   OR2_X1 i_0_0_0 (.A1(carryWires), .A2(n_0_16), .ZN(sum[32]));
   halfAdder__0_11 genblk1_0_HA (.in1(coutWire), .in2(n_0_0), .cout(n_0_17), 
      .sum(sum[16]));
   halfAdder__0_14 genblk1_1_HA2 (.in1(n_0_1), .in2(n_0_17), .cout(n_0_18), 
      .sum(sum[17]));
   halfAdder__0_17 genblk1_2_HA2 (.in1(n_0_2), .in2(n_0_18), .cout(n_0_19), 
      .sum(sum[18]));
   halfAdder__0_20 genblk1_3_HA2 (.in1(n_0_3), .in2(n_0_19), .cout(n_0_20), 
      .sum(sum[19]));
   halfAdder__0_23 genblk1_4_HA2 (.in1(n_0_4), .in2(n_0_20), .cout(n_0_21), 
      .sum(sum[20]));
   halfAdder__0_26 genblk1_5_HA2 (.in1(n_0_5), .in2(n_0_21), .cout(n_0_22), 
      .sum(sum[21]));
   halfAdder__0_29 genblk1_6_HA2 (.in1(n_0_6), .in2(n_0_22), .cout(n_0_23), 
      .sum(sum[22]));
   halfAdder__0_32 genblk1_7_HA2 (.in1(n_0_7), .in2(n_0_23), .cout(n_0_24), 
      .sum(sum[23]));
   halfAdder__0_35 genblk1_8_HA2 (.in1(n_0_8), .in2(n_0_24), .cout(n_0_25), 
      .sum(sum[24]));
   halfAdder__0_38 genblk1_9_HA2 (.in1(n_0_9), .in2(n_0_25), .cout(n_0_26), 
      .sum(sum[25]));
   halfAdder__0_41 genblk1_10_HA2 (.in1(n_0_10), .in2(n_0_26), .cout(n_0_27), 
      .sum(sum[26]));
   halfAdder__0_44 genblk1_11_HA2 (.in1(n_0_11), .in2(n_0_27), .cout(n_0_28), 
      .sum(sum[27]));
   halfAdder__0_47 genblk1_12_HA2 (.in1(n_0_12), .in2(n_0_28), .cout(n_0_29), 
      .sum(sum[28]));
   halfAdder__0_50 genblk1_13_HA2 (.in1(n_0_13), .in2(n_0_29), .cout(n_0_30), 
      .sum(sum[29]));
   halfAdder__0_53 genblk1_14_HA2 (.in1(n_0_14), .in2(n_0_30), .cout(n_0_31), 
      .sum(sum[30]));
   halfAdder genblk1_15_HA2 (.in1(n_0_15), .in2(n_0_31), .cout(carryWires), 
      .sum(sum[31]));
endmodule
