/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Nov  5 20:47:45 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2046132442 */

module n_case(A, B, S, enable);
   input [31:0]A;
   input [31:0]B;
   output [31:0]S;
   output enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;

   NOR4_X1 i_0_0 (.A1(n_0_60), .A2(n_0_57), .A3(n_0_43), .A4(n_0_0), .ZN(enable));
   NOR2_X1 i_0_1 (.A1(n_0_63), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   NOR4_X1 i_0_3 (.A1(B[29]), .A2(B[28]), .A3(B[27]), .A4(B[26]), .ZN(n_0_2));
   NOR4_X1 i_0_4 (.A1(B[30]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_3));
   AOI22_X1 i_0_5 (.A1(n_0_73), .A2(n_0_37), .B1(n_0_35), .B2(n_0_71), .ZN(S[0]));
   INV_X1 i_0_6 (.A(n_0_4), .ZN(S[1]));
   AOI22_X1 i_0_7 (.A1(A[1]), .A2(n_0_37), .B1(n_0_35), .B2(B[1]), .ZN(n_0_4));
   INV_X1 i_0_8 (.A(n_0_5), .ZN(S[2]));
   AOI22_X1 i_0_9 (.A1(A[2]), .A2(n_0_37), .B1(n_0_35), .B2(B[2]), .ZN(n_0_5));
   INV_X1 i_0_10 (.A(n_0_6), .ZN(S[3]));
   AOI22_X1 i_0_11 (.A1(A[3]), .A2(n_0_37), .B1(n_0_35), .B2(B[3]), .ZN(n_0_6));
   INV_X1 i_0_12 (.A(n_0_7), .ZN(S[4]));
   AOI22_X1 i_0_13 (.A1(A[4]), .A2(n_0_37), .B1(n_0_35), .B2(B[4]), .ZN(n_0_7));
   INV_X1 i_0_14 (.A(n_0_8), .ZN(S[5]));
   AOI22_X1 i_0_15 (.A1(A[5]), .A2(n_0_37), .B1(n_0_35), .B2(B[5]), .ZN(n_0_8));
   INV_X1 i_0_16 (.A(n_0_9), .ZN(S[6]));
   AOI22_X1 i_0_17 (.A1(A[6]), .A2(n_0_37), .B1(n_0_35), .B2(B[6]), .ZN(n_0_9));
   INV_X1 i_0_18 (.A(n_0_10), .ZN(S[7]));
   AOI22_X1 i_0_19 (.A1(A[7]), .A2(n_0_37), .B1(n_0_35), .B2(B[7]), .ZN(n_0_10));
   INV_X1 i_0_20 (.A(n_0_11), .ZN(S[8]));
   AOI22_X1 i_0_21 (.A1(A[8]), .A2(n_0_37), .B1(n_0_35), .B2(B[8]), .ZN(n_0_11));
   INV_X1 i_0_22 (.A(n_0_12), .ZN(S[9]));
   AOI22_X1 i_0_23 (.A1(A[9]), .A2(n_0_37), .B1(n_0_35), .B2(B[9]), .ZN(n_0_12));
   INV_X1 i_0_24 (.A(n_0_13), .ZN(S[10]));
   AOI22_X1 i_0_25 (.A1(A[10]), .A2(n_0_37), .B1(n_0_35), .B2(B[10]), .ZN(n_0_13));
   INV_X1 i_0_26 (.A(n_0_14), .ZN(S[11]));
   AOI22_X1 i_0_27 (.A1(A[11]), .A2(n_0_37), .B1(n_0_35), .B2(B[11]), .ZN(n_0_14));
   INV_X1 i_0_28 (.A(n_0_15), .ZN(S[12]));
   AOI22_X1 i_0_29 (.A1(A[12]), .A2(n_0_37), .B1(n_0_35), .B2(B[12]), .ZN(n_0_15));
   INV_X1 i_0_30 (.A(n_0_16), .ZN(S[13]));
   AOI22_X1 i_0_31 (.A1(A[13]), .A2(n_0_37), .B1(n_0_35), .B2(B[13]), .ZN(n_0_16));
   INV_X1 i_0_32 (.A(n_0_17), .ZN(S[14]));
   AOI22_X1 i_0_33 (.A1(A[14]), .A2(n_0_37), .B1(n_0_35), .B2(B[14]), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(n_0_18), .ZN(S[15]));
   AOI22_X1 i_0_35 (.A1(A[15]), .A2(n_0_37), .B1(n_0_35), .B2(B[15]), .ZN(n_0_18));
   INV_X1 i_0_36 (.A(n_0_19), .ZN(S[16]));
   AOI22_X1 i_0_37 (.A1(A[16]), .A2(n_0_37), .B1(n_0_35), .B2(B[16]), .ZN(n_0_19));
   INV_X1 i_0_38 (.A(n_0_20), .ZN(S[17]));
   AOI22_X1 i_0_39 (.A1(A[17]), .A2(n_0_37), .B1(n_0_35), .B2(B[17]), .ZN(n_0_20));
   INV_X1 i_0_40 (.A(n_0_21), .ZN(S[18]));
   AOI22_X1 i_0_41 (.A1(A[18]), .A2(n_0_37), .B1(n_0_35), .B2(B[18]), .ZN(n_0_21));
   INV_X1 i_0_42 (.A(n_0_22), .ZN(S[19]));
   AOI22_X1 i_0_43 (.A1(A[19]), .A2(n_0_37), .B1(n_0_35), .B2(B[19]), .ZN(n_0_22));
   INV_X1 i_0_44 (.A(n_0_23), .ZN(S[20]));
   AOI22_X1 i_0_45 (.A1(A[20]), .A2(n_0_37), .B1(n_0_35), .B2(B[20]), .ZN(n_0_23));
   INV_X1 i_0_46 (.A(n_0_24), .ZN(S[21]));
   AOI22_X1 i_0_47 (.A1(A[21]), .A2(n_0_37), .B1(n_0_35), .B2(B[21]), .ZN(n_0_24));
   INV_X1 i_0_48 (.A(n_0_25), .ZN(S[22]));
   AOI22_X1 i_0_49 (.A1(A[22]), .A2(n_0_37), .B1(n_0_35), .B2(B[22]), .ZN(n_0_25));
   INV_X1 i_0_50 (.A(n_0_26), .ZN(S[23]));
   OAI22_X1 i_0_51 (.A1(n_0_34), .A2(A[23]), .B1(B[23]), .B2(n_0_38), .ZN(n_0_26));
   INV_X1 i_0_52 (.A(n_0_27), .ZN(S[24]));
   OAI22_X1 i_0_53 (.A1(n_0_34), .A2(A[24]), .B1(B[24]), .B2(n_0_38), .ZN(n_0_27));
   INV_X1 i_0_54 (.A(n_0_28), .ZN(S[25]));
   OAI22_X1 i_0_55 (.A1(n_0_34), .A2(A[25]), .B1(B[25]), .B2(n_0_38), .ZN(n_0_28));
   INV_X1 i_0_56 (.A(n_0_29), .ZN(S[26]));
   OAI22_X1 i_0_57 (.A1(n_0_34), .A2(A[26]), .B1(B[26]), .B2(n_0_38), .ZN(n_0_29));
   INV_X1 i_0_58 (.A(n_0_30), .ZN(S[27]));
   OAI22_X1 i_0_59 (.A1(n_0_34), .A2(A[27]), .B1(B[27]), .B2(n_0_38), .ZN(n_0_30));
   INV_X1 i_0_60 (.A(n_0_31), .ZN(S[28]));
   OAI22_X1 i_0_61 (.A1(n_0_34), .A2(A[28]), .B1(B[28]), .B2(n_0_38), .ZN(n_0_31));
   INV_X1 i_0_62 (.A(n_0_32), .ZN(S[29]));
   OAI22_X1 i_0_63 (.A1(n_0_34), .A2(A[29]), .B1(B[29]), .B2(n_0_38), .ZN(n_0_32));
   INV_X1 i_0_64 (.A(n_0_33), .ZN(S[30]));
   OAI22_X1 i_0_65 (.A1(n_0_34), .A2(A[30]), .B1(B[30]), .B2(n_0_38), .ZN(n_0_33));
   OAI211_X1 i_0_66 (.A(n_0_48), .B(n_0_38), .C1(n_0_40), .C2(n_0_42), .ZN(
      n_0_34));
   AOI22_X1 i_0_67 (.A1(n_0_74), .A2(n_0_37), .B1(n_0_35), .B2(n_0_72), .ZN(
      S[31]));
   NOR2_X1 i_0_68 (.A1(n_0_36), .A2(n_0_38), .ZN(n_0_35));
   OAI21_X1 i_0_69 (.A(n_0_48), .B1(n_0_42), .B2(n_0_40), .ZN(n_0_36));
   AND3_X1 i_0_70 (.A1(n_0_48), .A2(n_0_38), .A3(n_0_39), .ZN(n_0_37));
   NOR2_X1 i_0_71 (.A1(n_0_47), .A2(n_0_43), .ZN(n_0_38));
   NAND2_X1 i_0_72 (.A1(n_0_41), .A2(n_0_42), .ZN(n_0_39));
   INV_X1 i_0_73 (.A(n_0_41), .ZN(n_0_40));
   AND2_X1 i_0_74 (.A1(n_0_60), .A2(n_0_57), .ZN(n_0_41));
   XNOR2_X1 i_0_75 (.A(n_0_74), .B(B[31]), .ZN(n_0_42));
   NOR2_X1 i_0_76 (.A1(n_0_49), .A2(n_0_44), .ZN(n_0_43));
   NAND2_X1 i_0_77 (.A1(n_0_46), .A2(n_0_45), .ZN(n_0_44));
   NOR4_X1 i_0_78 (.A1(A[29]), .A2(A[28]), .A3(A[27]), .A4(A[26]), .ZN(n_0_45));
   NOR4_X1 i_0_79 (.A1(A[30]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_46));
   NOR4_X1 i_0_80 (.A1(n_0_63), .A2(n_0_62), .A3(n_0_61), .A4(n_0_57), .ZN(
      n_0_47));
   AOI22_X1 i_0_81 (.A1(n_0_57), .A2(n_0_49), .B1(n_0_63), .B2(n_0_60), .ZN(
      n_0_48));
   NAND3_X1 i_0_82 (.A1(n_0_56), .A2(n_0_55), .A3(n_0_50), .ZN(n_0_49));
   AND4_X1 i_0_83 (.A1(n_0_54), .A2(n_0_53), .A3(n_0_52), .A4(n_0_51), .ZN(
      n_0_50));
   NOR3_X1 i_0_84 (.A1(A[10]), .A2(A[9]), .A3(A[8]), .ZN(n_0_51));
   NOR4_X1 i_0_85 (.A1(A[11]), .A2(A[7]), .A3(A[6]), .A4(A[4]), .ZN(n_0_52));
   NOR4_X1 i_0_86 (.A1(A[5]), .A2(A[3]), .A3(A[2]), .A4(A[1]), .ZN(n_0_53));
   NOR4_X1 i_0_87 (.A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[0]), .ZN(n_0_54));
   NOR4_X1 i_0_88 (.A1(A[19]), .A2(A[18]), .A3(A[16]), .A4(A[12]), .ZN(n_0_55));
   NOR4_X1 i_0_89 (.A1(A[17]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n_0_56));
   NOR2_X1 i_0_90 (.A1(n_0_59), .A2(n_0_58), .ZN(n_0_57));
   NAND4_X1 i_0_91 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_0_58));
   NAND4_X1 i_0_92 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_59));
   NOR2_X1 i_0_93 (.A1(n_0_62), .A2(n_0_61), .ZN(n_0_60));
   NAND4_X1 i_0_94 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_61));
   NAND4_X1 i_0_95 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_62));
   NAND3_X1 i_0_96 (.A1(n_0_66), .A2(n_0_65), .A3(n_0_64), .ZN(n_0_63));
   NOR4_X1 i_0_97 (.A1(B[19]), .A2(B[18]), .A3(B[16]), .A4(B[12]), .ZN(n_0_64));
   NOR4_X1 i_0_98 (.A1(B[17]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n_0_65));
   AND4_X1 i_0_99 (.A1(n_0_70), .A2(n_0_69), .A3(n_0_68), .A4(n_0_67), .ZN(
      n_0_66));
   NOR3_X1 i_0_100 (.A1(B[10]), .A2(B[9]), .A3(B[8]), .ZN(n_0_67));
   NOR4_X1 i_0_101 (.A1(B[11]), .A2(B[7]), .A3(B[6]), .A4(B[4]), .ZN(n_0_68));
   NOR4_X1 i_0_102 (.A1(B[5]), .A2(B[3]), .A3(B[2]), .A4(B[1]), .ZN(n_0_69));
   NOR4_X1 i_0_103 (.A1(B[22]), .A2(B[21]), .A3(B[20]), .A4(B[0]), .ZN(n_0_70));
   INV_X1 i_0_104 (.A(B[0]), .ZN(n_0_71));
   INV_X1 i_0_105 (.A(B[31]), .ZN(n_0_72));
   INV_X1 i_0_106 (.A(A[0]), .ZN(n_0_73));
   INV_X1 i_0_107 (.A(A[31]), .ZN(n_0_74));
endmodule

module selector(A, B, edata, NA, NB);
   input [31:0]A;
   input [31:0]B;
   output [1:0]edata;
   output [36:0]NA;
   output [36:0]NB;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   AND2_X1 i_0_0 (.A1(NB[27]), .A2(NA[27]), .ZN(edata[0]));
   XOR2_X1 i_0_1 (.A(NB[27]), .B(NA[27]), .Z(edata[1]));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .ZN(NA[27]));
   NOR4_X1 i_0_3 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_0_0));
   NOR4_X1 i_0_4 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(NB[27]));
   NOR4_X1 i_0_6 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_2));
   NOR4_X1 i_0_7 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_3));
endmodule

module n_subn(A, B, Comp, SA, SB, EO, MA, MB);
   input [36:0]A;
   input [36:0]B;
   output Comp;
   output SA;
   output SB;
   output [7:0]EO;
   output [27:0]MA;
   output [27:0]MB;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;

   INV_X1 i_0_0 (.A(A[4]), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(A[5]), .ZN(n_0_1));
   OAI211_X1 i_0_2 (.A(n_0_0), .B(B[4]), .C1(n_0_1), .C2(B[5]), .ZN(n_0_2));
   INV_X1 i_0_3 (.A(B[6]), .ZN(n_0_3));
   INV_X1 i_0_4 (.A(B[5]), .ZN(n_0_4));
   OAI221_X1 i_0_5 (.A(n_0_2), .B1(n_0_3), .B2(A[6]), .C1(A[5]), .C2(n_0_4), 
      .ZN(n_0_5));
   INV_X1 i_0_6 (.A(A[6]), .ZN(n_0_6));
   INV_X1 i_0_7 (.A(A[7]), .ZN(n_0_7));
   OAI221_X1 i_0_8 (.A(n_0_5), .B1(B[6]), .B2(n_0_6), .C1(n_0_7), .C2(B[7]), 
      .ZN(n_0_8));
   INV_X1 i_0_9 (.A(B[8]), .ZN(n_0_9));
   INV_X1 i_0_10 (.A(B[7]), .ZN(n_0_10));
   OAI221_X1 i_0_11 (.A(n_0_8), .B1(n_0_9), .B2(A[8]), .C1(A[7]), .C2(n_0_10), 
      .ZN(n_0_11));
   INV_X1 i_0_12 (.A(A[8]), .ZN(n_0_12));
   INV_X1 i_0_13 (.A(A[9]), .ZN(n_0_13));
   OAI221_X1 i_0_14 (.A(n_0_11), .B1(B[8]), .B2(n_0_12), .C1(n_0_13), .C2(B[9]), 
      .ZN(n_0_14));
   INV_X1 i_0_15 (.A(B[10]), .ZN(n_0_15));
   INV_X1 i_0_16 (.A(B[9]), .ZN(n_0_16));
   OAI221_X1 i_0_17 (.A(n_0_14), .B1(n_0_15), .B2(A[10]), .C1(A[9]), .C2(n_0_16), 
      .ZN(n_0_17));
   INV_X1 i_0_18 (.A(A[10]), .ZN(n_0_18));
   INV_X1 i_0_19 (.A(A[11]), .ZN(n_0_19));
   OAI221_X1 i_0_20 (.A(n_0_17), .B1(B[10]), .B2(n_0_18), .C1(n_0_19), .C2(B[11]), 
      .ZN(n_0_20));
   INV_X1 i_0_21 (.A(B[12]), .ZN(n_0_21));
   INV_X1 i_0_22 (.A(B[11]), .ZN(n_0_22));
   OAI221_X1 i_0_23 (.A(n_0_20), .B1(n_0_21), .B2(A[12]), .C1(A[11]), .C2(n_0_22), 
      .ZN(n_0_23));
   INV_X1 i_0_24 (.A(A[12]), .ZN(n_0_24));
   INV_X1 i_0_25 (.A(A[13]), .ZN(n_0_25));
   OAI221_X1 i_0_26 (.A(n_0_23), .B1(B[12]), .B2(n_0_24), .C1(n_0_25), .C2(B[13]), 
      .ZN(n_0_26));
   INV_X1 i_0_27 (.A(B[14]), .ZN(n_0_27));
   INV_X1 i_0_28 (.A(B[13]), .ZN(n_0_28));
   OAI221_X1 i_0_29 (.A(n_0_26), .B1(n_0_27), .B2(A[14]), .C1(A[13]), .C2(n_0_28), 
      .ZN(n_0_29));
   INV_X1 i_0_30 (.A(A[14]), .ZN(n_0_30));
   INV_X1 i_0_31 (.A(A[15]), .ZN(n_0_31));
   OAI221_X1 i_0_32 (.A(n_0_29), .B1(B[14]), .B2(n_0_30), .C1(n_0_31), .C2(B[15]), 
      .ZN(n_0_32));
   INV_X1 i_0_33 (.A(B[15]), .ZN(n_0_33));
   INV_X1 i_0_34 (.A(B[16]), .ZN(n_0_34));
   OAI221_X1 i_0_35 (.A(n_0_32), .B1(A[15]), .B2(n_0_33), .C1(n_0_34), .C2(A[16]), 
      .ZN(n_0_35));
   INV_X1 i_0_36 (.A(B[17]), .ZN(n_0_36));
   AOI22_X1 i_0_37 (.A1(n_0_34), .A2(A[16]), .B1(n_0_36), .B2(A[17]), .ZN(n_0_37));
   INV_X1 i_0_38 (.A(A[17]), .ZN(n_0_38));
   AOI22_X1 i_0_39 (.A1(n_0_35), .A2(n_0_37), .B1(n_0_38), .B2(B[17]), .ZN(
      n_0_39));
   INV_X1 i_0_40 (.A(B[18]), .ZN(n_0_40));
   AOI21_X1 i_0_41 (.A(n_0_39), .B1(A[18]), .B2(n_0_40), .ZN(n_0_41));
   INV_X1 i_0_42 (.A(A[18]), .ZN(n_0_42));
   INV_X1 i_0_43 (.A(A[19]), .ZN(n_0_43));
   AOI221_X1 i_0_44 (.A(n_0_41), .B1(n_0_42), .B2(B[18]), .C1(B[19]), .C2(n_0_43), 
      .ZN(n_0_44));
   INV_X1 i_0_45 (.A(B[19]), .ZN(n_0_45));
   INV_X1 i_0_46 (.A(B[20]), .ZN(n_0_46));
   AOI221_X1 i_0_47 (.A(n_0_44), .B1(n_0_45), .B2(A[19]), .C1(A[20]), .C2(n_0_46), 
      .ZN(n_0_47));
   INV_X1 i_0_48 (.A(A[20]), .ZN(n_0_48));
   INV_X1 i_0_49 (.A(A[21]), .ZN(n_0_49));
   AOI221_X1 i_0_50 (.A(n_0_47), .B1(n_0_48), .B2(B[20]), .C1(B[21]), .C2(n_0_49), 
      .ZN(n_0_50));
   INV_X1 i_0_51 (.A(B[21]), .ZN(n_0_51));
   INV_X1 i_0_52 (.A(B[22]), .ZN(n_0_52));
   AOI221_X1 i_0_53 (.A(n_0_50), .B1(n_0_51), .B2(A[21]), .C1(A[22]), .C2(n_0_52), 
      .ZN(n_0_53));
   INV_X1 i_0_54 (.A(A[22]), .ZN(n_0_54));
   INV_X1 i_0_55 (.A(A[23]), .ZN(n_0_55));
   AOI221_X1 i_0_56 (.A(n_0_53), .B1(n_0_54), .B2(B[22]), .C1(B[23]), .C2(n_0_55), 
      .ZN(n_0_56));
   INV_X1 i_0_57 (.A(B[23]), .ZN(n_0_57));
   INV_X1 i_0_58 (.A(B[24]), .ZN(n_0_58));
   AOI221_X1 i_0_59 (.A(n_0_56), .B1(n_0_57), .B2(A[23]), .C1(A[24]), .C2(n_0_58), 
      .ZN(n_0_59));
   INV_X1 i_0_60 (.A(A[24]), .ZN(n_0_60));
   INV_X1 i_0_61 (.A(A[25]), .ZN(n_0_61));
   AOI221_X1 i_0_62 (.A(n_0_59), .B1(n_0_60), .B2(B[24]), .C1(B[25]), .C2(n_0_61), 
      .ZN(n_0_62));
   INV_X1 i_0_63 (.A(B[26]), .ZN(n_0_63));
   INV_X1 i_0_64 (.A(B[25]), .ZN(n_0_64));
   AOI221_X1 i_0_65 (.A(n_0_62), .B1(A[26]), .B2(n_0_63), .C1(n_0_64), .C2(A[25]), 
      .ZN(n_0_65));
   INV_X1 i_0_66 (.A(B[27]), .ZN(n_0_66));
   OAI22_X1 i_0_67 (.A1(n_0_63), .A2(A[26]), .B1(n_0_66), .B2(A[27]), .ZN(n_0_67));
   INV_X1 i_0_68 (.A(A[27]), .ZN(n_0_68));
   OAI22_X1 i_0_69 (.A1(n_0_65), .A2(n_0_67), .B1(B[27]), .B2(n_0_68), .ZN(Comp));
   INV_X1 i_0_70 (.A(Comp), .ZN(n_0_69));
   INV_X1 i_0_71 (.A(B[4]), .ZN(n_0_70));
   OAI22_X1 i_0_72 (.A1(n_0_69), .A2(n_0_70), .B1(Comp), .B2(n_0_0), .ZN(MB[4]));
   OAI22_X1 i_0_73 (.A1(n_0_69), .A2(n_0_4), .B1(n_0_1), .B2(Comp), .ZN(MB[5]));
   AOI22_X1 i_0_74 (.A1(n_0_69), .A2(n_0_6), .B1(n_0_3), .B2(Comp), .ZN(MB[6]));
   AOI22_X1 i_0_75 (.A1(n_0_69), .A2(n_0_7), .B1(n_0_10), .B2(Comp), .ZN(MB[7]));
   AOI22_X1 i_0_76 (.A1(n_0_69), .A2(n_0_12), .B1(n_0_9), .B2(Comp), .ZN(MB[8]));
   AOI22_X1 i_0_77 (.A1(n_0_69), .A2(n_0_13), .B1(n_0_16), .B2(Comp), .ZN(MB[9]));
   AOI22_X1 i_0_78 (.A1(n_0_69), .A2(n_0_18), .B1(n_0_15), .B2(Comp), .ZN(MB[10]));
   AOI22_X1 i_0_79 (.A1(n_0_69), .A2(n_0_19), .B1(n_0_22), .B2(Comp), .ZN(MB[11]));
   AOI22_X1 i_0_80 (.A1(n_0_69), .A2(n_0_24), .B1(n_0_21), .B2(Comp), .ZN(MB[12]));
   AOI22_X1 i_0_81 (.A1(n_0_69), .A2(n_0_25), .B1(n_0_28), .B2(Comp), .ZN(MB[13]));
   AOI22_X1 i_0_82 (.A1(n_0_69), .A2(n_0_30), .B1(n_0_27), .B2(Comp), .ZN(MB[14]));
   AOI22_X1 i_0_83 (.A1(n_0_69), .A2(n_0_31), .B1(n_0_33), .B2(Comp), .ZN(MB[15]));
   INV_X1 i_0_84 (.A(A[16]), .ZN(n_0_71));
   AOI22_X1 i_0_85 (.A1(n_0_69), .A2(n_0_71), .B1(n_0_34), .B2(Comp), .ZN(MB[16]));
   AOI22_X1 i_0_86 (.A1(n_0_69), .A2(n_0_38), .B1(n_0_36), .B2(Comp), .ZN(MB[17]));
   OAI22_X1 i_0_87 (.A1(n_0_69), .A2(n_0_40), .B1(n_0_42), .B2(Comp), .ZN(MB[18]));
   AOI22_X1 i_0_88 (.A1(n_0_69), .A2(n_0_43), .B1(n_0_45), .B2(Comp), .ZN(MB[19]));
   OAI22_X1 i_0_89 (.A1(n_0_69), .A2(n_0_46), .B1(n_0_48), .B2(Comp), .ZN(MB[20]));
   AOI22_X1 i_0_90 (.A1(n_0_69), .A2(n_0_49), .B1(n_0_51), .B2(Comp), .ZN(MB[21]));
   OAI22_X1 i_0_91 (.A1(n_0_69), .A2(n_0_52), .B1(n_0_54), .B2(Comp), .ZN(MB[22]));
   AOI22_X1 i_0_92 (.A1(n_0_69), .A2(n_0_55), .B1(n_0_57), .B2(Comp), .ZN(MB[23]));
   OAI22_X1 i_0_93 (.A1(n_0_69), .A2(n_0_58), .B1(n_0_60), .B2(Comp), .ZN(MB[24]));
   AOI22_X1 i_0_94 (.A1(n_0_69), .A2(n_0_61), .B1(n_0_64), .B2(Comp), .ZN(MB[25]));
   INV_X1 i_0_95 (.A(A[26]), .ZN(n_0_72));
   OAI22_X1 i_0_96 (.A1(n_0_69), .A2(n_0_63), .B1(n_0_72), .B2(Comp), .ZN(MB[26]));
   NOR2_X1 i_0_97 (.A1(n_0_66), .A2(n_0_68), .ZN(MB[27]));
   AOI22_X1 i_0_98 (.A1(n_0_69), .A2(n_0_70), .B1(Comp), .B2(n_0_0), .ZN(MA[4]));
   AOI22_X1 i_0_99 (.A1(n_0_69), .A2(n_0_4), .B1(n_0_1), .B2(Comp), .ZN(MA[5]));
   OAI22_X1 i_0_100 (.A1(n_0_69), .A2(n_0_6), .B1(n_0_3), .B2(Comp), .ZN(MA[6]));
   OAI22_X1 i_0_101 (.A1(n_0_69), .A2(n_0_7), .B1(n_0_10), .B2(Comp), .ZN(MA[7]));
   OAI22_X1 i_0_102 (.A1(n_0_69), .A2(n_0_12), .B1(n_0_9), .B2(Comp), .ZN(MA[8]));
   OAI22_X1 i_0_103 (.A1(n_0_69), .A2(n_0_13), .B1(n_0_16), .B2(Comp), .ZN(MA[9]));
   OAI22_X1 i_0_104 (.A1(n_0_69), .A2(n_0_18), .B1(n_0_15), .B2(Comp), .ZN(
      MA[10]));
   OAI22_X1 i_0_105 (.A1(n_0_69), .A2(n_0_19), .B1(n_0_22), .B2(Comp), .ZN(
      MA[11]));
   OAI22_X1 i_0_106 (.A1(n_0_69), .A2(n_0_24), .B1(n_0_21), .B2(Comp), .ZN(
      MA[12]));
   OAI22_X1 i_0_107 (.A1(n_0_69), .A2(n_0_25), .B1(n_0_28), .B2(Comp), .ZN(
      MA[13]));
   OAI22_X1 i_0_108 (.A1(n_0_69), .A2(n_0_30), .B1(n_0_27), .B2(Comp), .ZN(
      MA[14]));
   OAI22_X1 i_0_109 (.A1(n_0_69), .A2(n_0_31), .B1(n_0_33), .B2(Comp), .ZN(
      MA[15]));
   OAI22_X1 i_0_110 (.A1(n_0_69), .A2(n_0_71), .B1(n_0_34), .B2(Comp), .ZN(
      MA[16]));
   OAI22_X1 i_0_111 (.A1(n_0_69), .A2(n_0_38), .B1(n_0_36), .B2(Comp), .ZN(
      MA[17]));
   AOI22_X1 i_0_112 (.A1(n_0_69), .A2(n_0_40), .B1(n_0_42), .B2(Comp), .ZN(
      MA[18]));
   OAI22_X1 i_0_113 (.A1(n_0_69), .A2(n_0_43), .B1(n_0_45), .B2(Comp), .ZN(
      MA[19]));
   AOI22_X1 i_0_114 (.A1(n_0_69), .A2(n_0_46), .B1(n_0_48), .B2(Comp), .ZN(
      MA[20]));
   OAI22_X1 i_0_115 (.A1(n_0_69), .A2(n_0_49), .B1(n_0_51), .B2(Comp), .ZN(
      MA[21]));
   AOI22_X1 i_0_116 (.A1(n_0_69), .A2(n_0_52), .B1(n_0_54), .B2(Comp), .ZN(
      MA[22]));
   OAI22_X1 i_0_117 (.A1(n_0_69), .A2(n_0_55), .B1(n_0_57), .B2(Comp), .ZN(
      MA[23]));
   AOI22_X1 i_0_118 (.A1(n_0_69), .A2(n_0_58), .B1(n_0_60), .B2(Comp), .ZN(
      MA[24]));
   OAI22_X1 i_0_119 (.A1(n_0_69), .A2(n_0_61), .B1(n_0_64), .B2(Comp), .ZN(
      MA[25]));
   AOI22_X1 i_0_120 (.A1(n_0_69), .A2(n_0_63), .B1(n_0_72), .B2(Comp), .ZN(
      MA[26]));
   NAND2_X1 i_0_121 (.A1(n_0_66), .A2(n_0_68), .ZN(MA[27]));
endmodule

module comp_exp(A, B, edata, SA, SB, Comp, Enor, MMax, MShift, Dexp);
   input [36:0]A;
   input [36:0]B;
   input [1:0]edata;
   output SA;
   output SB;
   output Comp;
   output [7:0]Enor;
   output [27:0]MMax;
   output [27:0]MShift;
   output [4:0]Dexp;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(Dexp[0]));
   OAI211_X1 i_0_1 (.A(n_0_29), .B(n_0_2), .C1(n_0_31), .C2(n_0_30), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(Dexp[1]));
   OAI211_X1 i_0_3 (.A(n_0_27), .B(n_0_2), .C1(n_0_32), .C2(n_0_28), .ZN(n_0_1));
   AOI21_X1 i_0_4 (.A(n_0_8), .B1(n_0_6), .B2(n_0_3), .ZN(n_0_2));
   NOR2_X1 i_0_5 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(n_0_7), .A2(n_0_4), .ZN(Dexp[2]));
   XOR2_X1 i_0_7 (.A(n_0_26), .B(n_0_25), .Z(n_0_4));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_5), .ZN(Dexp[3]));
   XNOR2_X1 i_0_9 (.A(n_0_24), .B(n_0_23), .ZN(n_0_5));
   OR2_X1 i_0_10 (.A1(n_0_8), .A2(n_0_6), .ZN(Dexp[4]));
   XOR2_X1 i_0_11 (.A(n_0_21), .B(n_0_20), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   OAI22_X1 i_0_13 (.A1(n_0_34), .A2(n_0_13), .B1(n_0_16), .B2(n_0_9), .ZN(n_0_8));
   AOI211_X1 i_0_14 (.A(n_0_10), .B(n_0_19), .C1(n_0_65), .C2(n_0_11), .ZN(n_0_9));
   NOR2_X1 i_0_15 (.A1(n_0_64), .A2(n_0_11), .ZN(n_0_10));
   XOR2_X1 i_0_16 (.A(Comp), .B(n_0_12), .Z(n_0_11));
   NOR2_X1 i_0_17 (.A1(n_0_67), .A2(n_0_52), .ZN(n_0_12));
   NOR3_X1 i_0_18 (.A1(n_0_15), .A2(n_0_14), .A3(n_0_16), .ZN(n_0_13));
   OAI33_X1 i_0_19 (.A1(n_0_52), .A2(n_0_17), .A3(n_0_41), .B1(A[34]), .B2(
      n_0_65), .B3(Comp), .ZN(n_0_14));
   AOI211_X1 i_0_20 (.A(n_0_156), .B(Comp), .C1(A[34]), .C2(n_0_65), .ZN(n_0_15));
   NOR4_X1 i_0_21 (.A1(n_0_67), .A2(n_0_64), .A3(n_0_49), .A4(n_0_18), .ZN(
      n_0_16));
   NOR2_X1 i_0_22 (.A1(n_0_67), .A2(n_0_64), .ZN(n_0_17));
   INV_X1 i_0_23 (.A(n_0_19), .ZN(n_0_18));
   OAI21_X1 i_0_24 (.A(n_0_39), .B1(n_0_21), .B2(n_0_20), .ZN(n_0_19));
   OAI22_X1 i_0_25 (.A1(B[32]), .A2(n_0_123), .B1(n_0_154), .B2(A[32]), .ZN(
      n_0_20));
   INV_X1 i_0_26 (.A(n_0_22), .ZN(n_0_21));
   OAI21_X1 i_0_27 (.A(n_0_37), .B1(n_0_24), .B2(n_0_23), .ZN(n_0_22));
   OAI22_X1 i_0_28 (.A1(n_0_153), .A2(A[31]), .B1(B[31]), .B2(n_0_122), .ZN(
      n_0_23));
   OAI22_X1 i_0_29 (.A1(Enor[2]), .A2(n_0_33), .B1(n_0_26), .B2(n_0_25), 
      .ZN(n_0_24));
   OAI22_X1 i_0_30 (.A1(B[30]), .A2(n_0_121), .B1(n_0_152), .B2(A[30]), .ZN(
      n_0_25));
   NAND2_X1 i_0_31 (.A1(n_0_36), .A2(n_0_27), .ZN(n_0_26));
   NAND2_X1 i_0_32 (.A1(n_0_32), .A2(n_0_28), .ZN(n_0_27));
   OAI221_X1 i_0_33 (.A(n_0_29), .B1(n_0_47), .B2(n_0_41), .C1(A[28]), .C2(
      n_0_35), .ZN(n_0_28));
   NAND2_X1 i_0_34 (.A1(n_0_31), .A2(n_0_30), .ZN(n_0_29));
   NAND2_X1 i_0_35 (.A1(edata[1]), .A2(n_0_94), .ZN(n_0_30));
   AOI21_X1 i_0_36 (.A(n_0_48), .B1(B[28]), .B2(n_0_119), .ZN(n_0_31));
   NOR2_X1 i_0_37 (.A1(n_0_60), .A2(n_0_58), .ZN(n_0_32));
   NOR2_X1 i_0_38 (.A1(B[30]), .A2(A[30]), .ZN(n_0_33));
   AOI22_X1 i_0_39 (.A1(B[35]), .A2(n_0_126), .B1(n_0_157), .B2(A[35]), .ZN(
      n_0_34));
   OAI22_X1 i_0_40 (.A1(n_0_127), .A2(n_0_41), .B1(n_0_95), .B2(Comp), .ZN(
      MShift[4]));
   OAI22_X1 i_0_41 (.A1(n_0_128), .A2(n_0_41), .B1(n_0_96), .B2(Comp), .ZN(
      MShift[5]));
   OAI22_X1 i_0_42 (.A1(n_0_129), .A2(n_0_41), .B1(n_0_97), .B2(Comp), .ZN(
      MShift[6]));
   OAI22_X1 i_0_43 (.A1(n_0_130), .A2(n_0_41), .B1(n_0_98), .B2(Comp), .ZN(
      MShift[7]));
   OAI22_X1 i_0_44 (.A1(n_0_131), .A2(n_0_41), .B1(n_0_99), .B2(Comp), .ZN(
      MShift[8]));
   OAI22_X1 i_0_45 (.A1(n_0_132), .A2(n_0_41), .B1(n_0_100), .B2(Comp), .ZN(
      MShift[9]));
   OAI22_X1 i_0_46 (.A1(n_0_133), .A2(n_0_41), .B1(n_0_101), .B2(Comp), .ZN(
      MShift[10]));
   OAI22_X1 i_0_47 (.A1(n_0_134), .A2(n_0_41), .B1(n_0_102), .B2(Comp), .ZN(
      MShift[11]));
   OAI22_X1 i_0_48 (.A1(n_0_135), .A2(n_0_41), .B1(n_0_103), .B2(Comp), .ZN(
      MShift[12]));
   OAI22_X1 i_0_49 (.A1(n_0_136), .A2(n_0_41), .B1(n_0_104), .B2(Comp), .ZN(
      MShift[13]));
   OAI22_X1 i_0_50 (.A1(n_0_137), .A2(n_0_41), .B1(n_0_105), .B2(Comp), .ZN(
      MShift[14]));
   OAI22_X1 i_0_51 (.A1(n_0_138), .A2(n_0_41), .B1(n_0_106), .B2(Comp), .ZN(
      MShift[15]));
   OAI22_X1 i_0_52 (.A1(n_0_139), .A2(n_0_41), .B1(n_0_107), .B2(Comp), .ZN(
      MShift[16]));
   OAI22_X1 i_0_53 (.A1(n_0_140), .A2(n_0_41), .B1(n_0_108), .B2(Comp), .ZN(
      MShift[17]));
   OAI22_X1 i_0_54 (.A1(n_0_141), .A2(n_0_41), .B1(n_0_109), .B2(Comp), .ZN(
      MShift[18]));
   OAI22_X1 i_0_55 (.A1(n_0_142), .A2(n_0_41), .B1(n_0_110), .B2(Comp), .ZN(
      MShift[19]));
   OAI22_X1 i_0_56 (.A1(n_0_143), .A2(n_0_41), .B1(n_0_111), .B2(Comp), .ZN(
      MShift[20]));
   OAI22_X1 i_0_57 (.A1(n_0_144), .A2(n_0_41), .B1(n_0_112), .B2(Comp), .ZN(
      MShift[21]));
   OAI22_X1 i_0_58 (.A1(n_0_145), .A2(n_0_41), .B1(n_0_113), .B2(Comp), .ZN(
      MShift[22]));
   OAI22_X1 i_0_59 (.A1(n_0_146), .A2(n_0_41), .B1(n_0_114), .B2(Comp), .ZN(
      MShift[23]));
   OAI22_X1 i_0_60 (.A1(n_0_147), .A2(n_0_41), .B1(n_0_115), .B2(Comp), .ZN(
      MShift[24]));
   OAI22_X1 i_0_61 (.A1(n_0_148), .A2(n_0_41), .B1(n_0_116), .B2(Comp), .ZN(
      MShift[25]));
   OAI22_X1 i_0_62 (.A1(n_0_149), .A2(n_0_41), .B1(n_0_117), .B2(Comp), .ZN(
      MShift[26]));
   OAI22_X1 i_0_63 (.A1(n_0_150), .A2(n_0_41), .B1(n_0_118), .B2(Comp), .ZN(
      MShift[27]));
   OAI22_X1 i_0_64 (.A1(n_0_95), .A2(n_0_41), .B1(n_0_127), .B2(Comp), .ZN(
      MMax[4]));
   OAI22_X1 i_0_65 (.A1(n_0_96), .A2(n_0_41), .B1(n_0_128), .B2(Comp), .ZN(
      MMax[5]));
   OAI22_X1 i_0_66 (.A1(n_0_97), .A2(n_0_41), .B1(n_0_129), .B2(Comp), .ZN(
      MMax[6]));
   OAI22_X1 i_0_67 (.A1(n_0_98), .A2(n_0_41), .B1(n_0_130), .B2(Comp), .ZN(
      MMax[7]));
   OAI22_X1 i_0_68 (.A1(n_0_99), .A2(n_0_41), .B1(n_0_131), .B2(Comp), .ZN(
      MMax[8]));
   OAI22_X1 i_0_69 (.A1(n_0_100), .A2(n_0_41), .B1(n_0_132), .B2(Comp), .ZN(
      MMax[9]));
   OAI22_X1 i_0_70 (.A1(n_0_101), .A2(n_0_41), .B1(n_0_133), .B2(Comp), .ZN(
      MMax[10]));
   OAI22_X1 i_0_71 (.A1(n_0_102), .A2(n_0_41), .B1(n_0_134), .B2(Comp), .ZN(
      MMax[11]));
   OAI22_X1 i_0_72 (.A1(n_0_103), .A2(n_0_41), .B1(n_0_135), .B2(Comp), .ZN(
      MMax[12]));
   OAI22_X1 i_0_73 (.A1(n_0_104), .A2(n_0_41), .B1(n_0_136), .B2(Comp), .ZN(
      MMax[13]));
   OAI22_X1 i_0_74 (.A1(n_0_105), .A2(n_0_41), .B1(n_0_137), .B2(Comp), .ZN(
      MMax[14]));
   OAI22_X1 i_0_75 (.A1(n_0_106), .A2(n_0_41), .B1(n_0_138), .B2(Comp), .ZN(
      MMax[15]));
   OAI22_X1 i_0_76 (.A1(n_0_107), .A2(n_0_41), .B1(n_0_139), .B2(Comp), .ZN(
      MMax[16]));
   OAI22_X1 i_0_77 (.A1(n_0_108), .A2(n_0_41), .B1(n_0_140), .B2(Comp), .ZN(
      MMax[17]));
   OAI22_X1 i_0_78 (.A1(n_0_109), .A2(n_0_41), .B1(n_0_141), .B2(Comp), .ZN(
      MMax[18]));
   OAI22_X1 i_0_79 (.A1(n_0_110), .A2(n_0_41), .B1(n_0_142), .B2(Comp), .ZN(
      MMax[19]));
   OAI22_X1 i_0_80 (.A1(n_0_111), .A2(n_0_41), .B1(n_0_143), .B2(Comp), .ZN(
      MMax[20]));
   OAI22_X1 i_0_81 (.A1(n_0_112), .A2(n_0_41), .B1(n_0_144), .B2(Comp), .ZN(
      MMax[21]));
   OAI22_X1 i_0_82 (.A1(n_0_113), .A2(n_0_41), .B1(n_0_145), .B2(Comp), .ZN(
      MMax[22]));
   OAI22_X1 i_0_83 (.A1(n_0_114), .A2(n_0_41), .B1(n_0_146), .B2(Comp), .ZN(
      MMax[23]));
   OAI22_X1 i_0_84 (.A1(n_0_115), .A2(n_0_41), .B1(n_0_147), .B2(Comp), .ZN(
      MMax[24]));
   OAI22_X1 i_0_85 (.A1(n_0_116), .A2(n_0_41), .B1(n_0_148), .B2(Comp), .ZN(
      MMax[25]));
   OAI22_X1 i_0_86 (.A1(n_0_117), .A2(n_0_41), .B1(n_0_149), .B2(Comp), .ZN(
      MMax[26]));
   OAI22_X1 i_0_87 (.A1(n_0_118), .A2(n_0_41), .B1(n_0_150), .B2(Comp), .ZN(
      MMax[27]));
   OAI21_X1 i_0_88 (.A(n_0_35), .B1(n_0_119), .B2(n_0_41), .ZN(Enor[0]));
   NAND2_X1 i_0_89 (.A1(B[28]), .A2(n_0_41), .ZN(n_0_35));
   OAI21_X1 i_0_90 (.A(n_0_36), .B1(n_0_151), .B2(n_0_120), .ZN(Enor[1]));
   OAI22_X1 i_0_91 (.A1(n_0_60), .A2(Comp), .B1(n_0_58), .B2(n_0_41), .ZN(n_0_36));
   OAI22_X1 i_0_92 (.A1(n_0_121), .A2(n_0_41), .B1(n_0_152), .B2(Comp), .ZN(
      Enor[2]));
   OAI21_X1 i_0_93 (.A(n_0_37), .B1(n_0_153), .B2(n_0_122), .ZN(Enor[3]));
   INV_X1 i_0_94 (.A(n_0_38), .ZN(n_0_37));
   OAI33_X1 i_0_95 (.A1(B[31]), .A2(n_0_122), .A3(n_0_41), .B1(n_0_153), 
      .B2(A[31]), .B3(Comp), .ZN(n_0_38));
   OAI21_X1 i_0_96 (.A(n_0_39), .B1(n_0_154), .B2(n_0_123), .ZN(Enor[4]));
   INV_X1 i_0_97 (.A(n_0_40), .ZN(n_0_39));
   OAI33_X1 i_0_98 (.A1(B[32]), .A2(n_0_123), .A3(n_0_41), .B1(n_0_154), 
      .B2(A[32]), .B3(Comp), .ZN(n_0_40));
   OAI22_X1 i_0_99 (.A1(n_0_124), .A2(n_0_41), .B1(n_0_155), .B2(Comp), .ZN(
      Enor[5]));
   OAI22_X1 i_0_100 (.A1(n_0_125), .A2(n_0_41), .B1(n_0_156), .B2(Comp), 
      .ZN(Enor[6]));
   INV_X1 i_0_101 (.A(Comp), .ZN(n_0_41));
   OAI211_X1 i_0_102 (.A(n_0_42), .B(n_0_50), .C1(B[35]), .C2(n_0_126), .ZN(Comp));
   OAI22_X1 i_0_103 (.A1(n_0_157), .A2(A[35]), .B1(n_0_67), .B2(n_0_43), 
      .ZN(n_0_42));
   AOI21_X1 i_0_104 (.A(n_0_49), .B1(n_0_63), .B2(n_0_44), .ZN(n_0_43));
   OAI21_X1 i_0_105 (.A(n_0_62), .B1(n_0_61), .B2(n_0_45), .ZN(n_0_44));
   INV_X1 i_0_106 (.A(n_0_46), .ZN(n_0_45));
   OAI21_X1 i_0_107 (.A(n_0_59), .B1(n_0_58), .B2(n_0_48), .ZN(n_0_46));
   INV_X1 i_0_108 (.A(n_0_48), .ZN(n_0_47));
   NOR2_X1 i_0_109 (.A1(B[28]), .A2(n_0_119), .ZN(n_0_48));
   OAI21_X1 i_0_110 (.A(n_0_65), .B1(n_0_156), .B2(A[34]), .ZN(n_0_49));
   OAI211_X1 i_0_111 (.A(n_0_51), .B(n_0_68), .C1(n_0_67), .C2(n_0_53), .ZN(
      n_0_50));
   AOI221_X1 i_0_112 (.A(n_0_52), .B1(B[35]), .B2(n_0_126), .C1(B[27]), .C2(
      n_0_118), .ZN(n_0_51));
   NOR2_X1 i_0_113 (.A1(n_0_156), .A2(A[34]), .ZN(n_0_52));
   AOI21_X1 i_0_114 (.A(n_0_66), .B1(n_0_63), .B2(n_0_54), .ZN(n_0_53));
   OAI21_X1 i_0_115 (.A(n_0_62), .B1(n_0_61), .B2(n_0_55), .ZN(n_0_54));
   INV_X1 i_0_116 (.A(n_0_56), .ZN(n_0_55));
   OAI21_X1 i_0_117 (.A(n_0_59), .B1(n_0_58), .B2(n_0_57), .ZN(n_0_56));
   NAND2_X1 i_0_118 (.A1(B[28]), .A2(n_0_119), .ZN(n_0_57));
   NOR2_X1 i_0_119 (.A1(B[29]), .A2(n_0_120), .ZN(n_0_58));
   AOI21_X1 i_0_120 (.A(n_0_60), .B1(B[30]), .B2(n_0_121), .ZN(n_0_59));
   NOR2_X1 i_0_121 (.A1(n_0_151), .A2(A[29]), .ZN(n_0_60));
   OAI22_X1 i_0_122 (.A1(B[31]), .A2(n_0_122), .B1(B[30]), .B2(n_0_121), 
      .ZN(n_0_61));
   AOI22_X1 i_0_123 (.A1(B[31]), .A2(n_0_122), .B1(B[32]), .B2(n_0_123), 
      .ZN(n_0_62));
   AOI21_X1 i_0_124 (.A(n_0_64), .B1(n_0_154), .B2(A[32]), .ZN(n_0_63));
   NOR2_X1 i_0_125 (.A1(B[33]), .A2(n_0_124), .ZN(n_0_64));
   INV_X1 i_0_126 (.A(n_0_66), .ZN(n_0_65));
   NOR2_X1 i_0_127 (.A1(n_0_155), .A2(A[33]), .ZN(n_0_66));
   NOR2_X1 i_0_128 (.A1(B[34]), .A2(n_0_125), .ZN(n_0_67));
   OAI221_X1 i_0_129 (.A(n_0_69), .B1(B[26]), .B2(n_0_117), .C1(B[27]), .C2(
      n_0_118), .ZN(n_0_68));
   OAI221_X1 i_0_130 (.A(n_0_70), .B1(n_0_149), .B2(A[26]), .C1(n_0_148), 
      .C2(A[25]), .ZN(n_0_69));
   OAI221_X1 i_0_131 (.A(n_0_71), .B1(B[24]), .B2(n_0_115), .C1(B[25]), .C2(
      n_0_116), .ZN(n_0_70));
   OAI21_X1 i_0_132 (.A(n_0_72), .B1(n_0_147), .B2(A[24]), .ZN(n_0_71));
   OAI21_X1 i_0_133 (.A(n_0_73), .B1(B[23]), .B2(n_0_114), .ZN(n_0_72));
   OAI221_X1 i_0_134 (.A(n_0_74), .B1(n_0_145), .B2(A[22]), .C1(n_0_146), 
      .C2(A[23]), .ZN(n_0_73));
   OAI221_X1 i_0_135 (.A(n_0_75), .B1(B[21]), .B2(n_0_112), .C1(B[22]), .C2(
      n_0_113), .ZN(n_0_74));
   OAI221_X1 i_0_136 (.A(n_0_76), .B1(n_0_143), .B2(A[20]), .C1(n_0_144), 
      .C2(A[21]), .ZN(n_0_75));
   OAI221_X1 i_0_137 (.A(n_0_77), .B1(B[19]), .B2(n_0_110), .C1(B[20]), .C2(
      n_0_111), .ZN(n_0_76));
   OAI221_X1 i_0_138 (.A(n_0_78), .B1(n_0_141), .B2(A[18]), .C1(n_0_142), 
      .C2(A[19]), .ZN(n_0_77));
   OAI221_X1 i_0_139 (.A(n_0_79), .B1(B[17]), .B2(n_0_108), .C1(B[18]), .C2(
      n_0_109), .ZN(n_0_78));
   OAI221_X1 i_0_140 (.A(n_0_80), .B1(n_0_139), .B2(A[16]), .C1(n_0_140), 
      .C2(A[17]), .ZN(n_0_79));
   OAI221_X1 i_0_141 (.A(n_0_81), .B1(B[15]), .B2(n_0_106), .C1(B[16]), .C2(
      n_0_107), .ZN(n_0_80));
   OAI221_X1 i_0_142 (.A(n_0_82), .B1(n_0_137), .B2(A[14]), .C1(n_0_138), 
      .C2(A[15]), .ZN(n_0_81));
   OAI221_X1 i_0_143 (.A(n_0_83), .B1(B[13]), .B2(n_0_104), .C1(B[14]), .C2(
      n_0_105), .ZN(n_0_82));
   OAI221_X1 i_0_144 (.A(n_0_84), .B1(n_0_135), .B2(A[12]), .C1(n_0_136), 
      .C2(A[13]), .ZN(n_0_83));
   OAI221_X1 i_0_145 (.A(n_0_85), .B1(B[11]), .B2(n_0_102), .C1(B[12]), .C2(
      n_0_103), .ZN(n_0_84));
   OAI221_X1 i_0_146 (.A(n_0_86), .B1(n_0_133), .B2(A[10]), .C1(n_0_134), 
      .C2(A[11]), .ZN(n_0_85));
   OAI221_X1 i_0_147 (.A(n_0_87), .B1(B[9]), .B2(n_0_100), .C1(B[10]), .C2(
      n_0_101), .ZN(n_0_86));
   OAI221_X1 i_0_148 (.A(n_0_88), .B1(n_0_132), .B2(A[9]), .C1(n_0_131), 
      .C2(A[8]), .ZN(n_0_87));
   OAI221_X1 i_0_149 (.A(n_0_89), .B1(B[8]), .B2(n_0_99), .C1(B[7]), .C2(n_0_98), 
      .ZN(n_0_88));
   OAI221_X1 i_0_150 (.A(n_0_90), .B1(A[6]), .B2(n_0_91), .C1(n_0_130), .C2(A[7]), 
      .ZN(n_0_89));
   OAI21_X1 i_0_151 (.A(B[6]), .B1(n_0_97), .B2(n_0_92), .ZN(n_0_90));
   INV_X1 i_0_152 (.A(n_0_92), .ZN(n_0_91));
   OAI21_X1 i_0_153 (.A(n_0_93), .B1(n_0_128), .B2(A[5]), .ZN(n_0_92));
   OAI211_X1 i_0_154 (.A(B[4]), .B(n_0_95), .C1(B[5]), .C2(n_0_96), .ZN(n_0_93));
   NAND2_X1 i_0_155 (.A1(n_0_157), .A2(n_0_126), .ZN(Enor[7]));
   INV_X1 i_0_156 (.A(edata[0]), .ZN(n_0_94));
   INV_X1 i_0_157 (.A(A[4]), .ZN(n_0_95));
   INV_X1 i_0_158 (.A(A[5]), .ZN(n_0_96));
   INV_X1 i_0_159 (.A(A[6]), .ZN(n_0_97));
   INV_X1 i_0_160 (.A(A[7]), .ZN(n_0_98));
   INV_X1 i_0_161 (.A(A[8]), .ZN(n_0_99));
   INV_X1 i_0_162 (.A(A[9]), .ZN(n_0_100));
   INV_X1 i_0_163 (.A(A[10]), .ZN(n_0_101));
   INV_X1 i_0_164 (.A(A[11]), .ZN(n_0_102));
   INV_X1 i_0_165 (.A(A[12]), .ZN(n_0_103));
   INV_X1 i_0_166 (.A(A[13]), .ZN(n_0_104));
   INV_X1 i_0_167 (.A(A[14]), .ZN(n_0_105));
   INV_X1 i_0_168 (.A(A[15]), .ZN(n_0_106));
   INV_X1 i_0_169 (.A(A[16]), .ZN(n_0_107));
   INV_X1 i_0_170 (.A(A[17]), .ZN(n_0_108));
   INV_X1 i_0_171 (.A(A[18]), .ZN(n_0_109));
   INV_X1 i_0_172 (.A(A[19]), .ZN(n_0_110));
   INV_X1 i_0_173 (.A(A[20]), .ZN(n_0_111));
   INV_X1 i_0_174 (.A(A[21]), .ZN(n_0_112));
   INV_X1 i_0_175 (.A(A[22]), .ZN(n_0_113));
   INV_X1 i_0_176 (.A(A[23]), .ZN(n_0_114));
   INV_X1 i_0_177 (.A(A[24]), .ZN(n_0_115));
   INV_X1 i_0_178 (.A(A[25]), .ZN(n_0_116));
   INV_X1 i_0_179 (.A(A[26]), .ZN(n_0_117));
   INV_X1 i_0_180 (.A(A[27]), .ZN(n_0_118));
   INV_X1 i_0_181 (.A(A[28]), .ZN(n_0_119));
   INV_X1 i_0_182 (.A(A[29]), .ZN(n_0_120));
   INV_X1 i_0_183 (.A(A[30]), .ZN(n_0_121));
   INV_X1 i_0_184 (.A(A[31]), .ZN(n_0_122));
   INV_X1 i_0_185 (.A(A[32]), .ZN(n_0_123));
   INV_X1 i_0_186 (.A(A[33]), .ZN(n_0_124));
   INV_X1 i_0_187 (.A(A[34]), .ZN(n_0_125));
   INV_X1 i_0_188 (.A(A[35]), .ZN(n_0_126));
   INV_X1 i_0_189 (.A(B[4]), .ZN(n_0_127));
   INV_X1 i_0_190 (.A(B[5]), .ZN(n_0_128));
   INV_X1 i_0_191 (.A(B[6]), .ZN(n_0_129));
   INV_X1 i_0_192 (.A(B[7]), .ZN(n_0_130));
   INV_X1 i_0_193 (.A(B[8]), .ZN(n_0_131));
   INV_X1 i_0_194 (.A(B[9]), .ZN(n_0_132));
   INV_X1 i_0_195 (.A(B[10]), .ZN(n_0_133));
   INV_X1 i_0_196 (.A(B[11]), .ZN(n_0_134));
   INV_X1 i_0_197 (.A(B[12]), .ZN(n_0_135));
   INV_X1 i_0_198 (.A(B[13]), .ZN(n_0_136));
   INV_X1 i_0_199 (.A(B[14]), .ZN(n_0_137));
   INV_X1 i_0_200 (.A(B[15]), .ZN(n_0_138));
   INV_X1 i_0_201 (.A(B[16]), .ZN(n_0_139));
   INV_X1 i_0_202 (.A(B[17]), .ZN(n_0_140));
   INV_X1 i_0_203 (.A(B[18]), .ZN(n_0_141));
   INV_X1 i_0_204 (.A(B[19]), .ZN(n_0_142));
   INV_X1 i_0_205 (.A(B[20]), .ZN(n_0_143));
   INV_X1 i_0_206 (.A(B[21]), .ZN(n_0_144));
   INV_X1 i_0_207 (.A(B[22]), .ZN(n_0_145));
   INV_X1 i_0_208 (.A(B[23]), .ZN(n_0_146));
   INV_X1 i_0_209 (.A(B[24]), .ZN(n_0_147));
   INV_X1 i_0_210 (.A(B[25]), .ZN(n_0_148));
   INV_X1 i_0_211 (.A(B[26]), .ZN(n_0_149));
   INV_X1 i_0_212 (.A(B[27]), .ZN(n_0_150));
   INV_X1 i_0_213 (.A(B[29]), .ZN(n_0_151));
   INV_X1 i_0_214 (.A(B[30]), .ZN(n_0_152));
   INV_X1 i_0_215 (.A(B[31]), .ZN(n_0_153));
   INV_X1 i_0_216 (.A(B[32]), .ZN(n_0_154));
   INV_X1 i_0_217 (.A(B[33]), .ZN(n_0_155));
   INV_X1 i_0_218 (.A(B[34]), .ZN(n_0_156));
   INV_X1 i_0_219 (.A(B[35]), .ZN(n_0_157));
endmodule

module mux2X1_r__0_355(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_357(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_359(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_361(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_363(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_365(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_367(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_369(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_371(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_373(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_375(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_377(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_379(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_381(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_383(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_385(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_387(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_389(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_391(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_393(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_395(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_397(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_399(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_401(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_403(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_405(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_407(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_409(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_411(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_413(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_415(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_417(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_419(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_421(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_423(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_425(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_427(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_429(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_431(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_433(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_435(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_437(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_439(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_441(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_443(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_445(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_447(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_449(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_451(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_453(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_455(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_457(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_459(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_461(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_463(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_465(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_467(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_469(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_471(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_473(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_475(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_477(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_479(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_481(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_483(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_485(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_487(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_489(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_491(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_493(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_495(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_497(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_499(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_501(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_503(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_505(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_507(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_509(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_511(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_513(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_515(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_517(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_519(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_521(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   AND2_X1 i_0_0 (.A1(sel), .A2(in0), .ZN(out));
endmodule

module mux2X1_r__0_523(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_525(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_527(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_529(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_531(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_533(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_535(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_537(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_539(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_541(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_543(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_545(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_547(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_549(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_551(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_553(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_555(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_557(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_559(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_561(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_563(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_565(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_567(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_569(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_571(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_573(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   AND2_X1 i_0_0 (.A1(sel), .A2(in0), .ZN(out));
endmodule

module mux2X1_r__0_575(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   AND2_X1 i_0_0 (.A1(sel), .A2(in0), .ZN(out));
endmodule

module mux2X1_r__0_579(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1_r__0_581(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_583(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_585(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_587(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_589(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_591(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_593(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_595(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_597(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_599(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_601(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_603(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_605(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_607(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_609(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_611(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_613(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_615(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_617(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_619(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_621(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_623(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_625(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1_r__0_627(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   AND2_X1 i_0_0 (.A1(sel), .A2(in0), .ZN(out));
endmodule

module n_shift_norm(shft, in, out);
   input [4:0]shft;
   input [27:0]in;
   output [27:0]out;

   wire [27:0]z4;
   wire [27:0]z3;
   wire [27:0]z2;
   wire [27:0]z1;

   mux2X1_r__0_355 genblk1_0_m9 (.in0(), .in1(z4[27]), .sel(shft[4]), .out(
      out[27]));
   mux2X1_r__0_357 genblk1_1_m9 (.in0(), .in1(z4[26]), .sel(shft[4]), .out(
      out[26]));
   mux2X1_r__0_359 genblk1_2_m9 (.in0(), .in1(z4[25]), .sel(shft[4]), .out(
      out[25]));
   mux2X1_r__0_361 genblk1_3_m9 (.in0(), .in1(z4[24]), .sel(shft[4]), .out(
      out[24]));
   mux2X1_r__0_363 genblk1_4_m9 (.in0(), .in1(z4[23]), .sel(shft[4]), .out(
      out[23]));
   mux2X1_r__0_365 genblk1_5_m9 (.in0(), .in1(z4[22]), .sel(shft[4]), .out(
      out[22]));
   mux2X1_r__0_367 genblk1_6_m9 (.in0(), .in1(z4[21]), .sel(shft[4]), .out(
      out[21]));
   mux2X1_r__0_369 genblk1_7_m9 (.in0(), .in1(z4[20]), .sel(shft[4]), .out(
      out[20]));
   mux2X1_r__0_371 genblk1_8_m9 (.in0(), .in1(z4[19]), .sel(shft[4]), .out(
      out[19]));
   mux2X1_r__0_373 genblk1_9_m9 (.in0(), .in1(z4[18]), .sel(shft[4]), .out(
      out[18]));
   mux2X1_r__0_375 genblk1_10_m9 (.in0(), .in1(z4[17]), .sel(shft[4]), .out(
      out[17]));
   mux2X1_r__0_377 genblk1_11_m9 (.in0(), .in1(z4[16]), .sel(shft[4]), .out(
      out[16]));
   mux2X1_r__0_379 genblk1_12_m9 (.in0(), .in1(z4[15]), .sel(shft[4]), .out(
      out[15]));
   mux2X1_r__0_381 genblk1_13_m9 (.in0(), .in1(z4[14]), .sel(shft[4]), .out(
      out[14]));
   mux2X1_r__0_383 genblk1_14_m9 (.in0(), .in1(z4[13]), .sel(shft[4]), .out(
      out[13]));
   mux2X1_r__0_385 genblk1_15_m9 (.in0(), .in1(z4[12]), .sel(shft[4]), .out(
      out[12]));
   mux2X1_r__0_387 genblk1_16_m10 (.in0(z4[27]), .in1(z4[11]), .sel(shft[4]), 
      .out(out[11]));
   mux2X1_r__0_389 genblk1_17_m10 (.in0(z4[26]), .in1(z4[10]), .sel(shft[4]), 
      .out(out[10]));
   mux2X1_r__0_391 genblk1_18_m10 (.in0(z4[25]), .in1(z4[9]), .sel(shft[4]), 
      .out(out[9]));
   mux2X1_r__0_393 genblk1_19_m10 (.in0(z4[24]), .in1(z4[8]), .sel(shft[4]), 
      .out(out[8]));
   mux2X1_r__0_395 genblk1_20_m10 (.in0(z4[23]), .in1(z4[7]), .sel(shft[4]), 
      .out(out[7]));
   mux2X1_r__0_397 genblk1_21_m10 (.in0(z4[22]), .in1(z4[6]), .sel(shft[4]), 
      .out(out[6]));
   mux2X1_r__0_399 genblk1_22_m10 (.in0(z4[21]), .in1(z4[5]), .sel(shft[4]), 
      .out(out[5]));
   mux2X1_r__0_401 genblk1_23_m10 (.in0(z4[20]), .in1(z4[4]), .sel(shft[4]), 
      .out(out[4]));
   mux2X1_r__0_403 genblk1_24_m10 (.in0(z4[19]), .in1(z4[3]), .sel(shft[4]), 
      .out(out[3]));
   mux2X1_r__0_405 genblk1_25_m10 (.in0(z4[18]), .in1(z4[2]), .sel(shft[4]), 
      .out(out[2]));
   mux2X1_r__0_407 genblk1_26_m10 (.in0(z4[17]), .in1(z4[1]), .sel(shft[4]), 
      .out(out[1]));
   mux2X1_r__0_409 genblk1_27_m10 (.in0(z4[16]), .in1(z4[0]), .sel(shft[4]), 
      .out(out[0]));
   mux2X1_r__0_411 genblk1_0_m7 (.in0(), .in1(z3[27]), .sel(shft[3]), .out(
      z4[27]));
   mux2X1_r__0_413 genblk1_1_m7 (.in0(), .in1(z3[26]), .sel(shft[3]), .out(
      z4[26]));
   mux2X1_r__0_415 genblk1_2_m7 (.in0(), .in1(z3[25]), .sel(shft[3]), .out(
      z4[25]));
   mux2X1_r__0_417 genblk1_3_m7 (.in0(), .in1(z3[24]), .sel(shft[3]), .out(
      z4[24]));
   mux2X1_r__0_419 genblk1_4_m7 (.in0(), .in1(z3[23]), .sel(shft[3]), .out(
      z4[23]));
   mux2X1_r__0_421 genblk1_5_m7 (.in0(), .in1(z3[22]), .sel(shft[3]), .out(
      z4[22]));
   mux2X1_r__0_423 genblk1_6_m7 (.in0(), .in1(z3[21]), .sel(shft[3]), .out(
      z4[21]));
   mux2X1_r__0_425 genblk1_7_m7 (.in0(), .in1(z3[20]), .sel(shft[3]), .out(
      z4[20]));
   mux2X1_r__0_427 genblk1_8_m8 (.in0(z3[27]), .in1(z3[19]), .sel(shft[3]), 
      .out(z4[19]));
   mux2X1_r__0_429 genblk1_9_m8 (.in0(z3[26]), .in1(z3[18]), .sel(shft[3]), 
      .out(z4[18]));
   mux2X1_r__0_431 genblk1_10_m8 (.in0(z3[25]), .in1(z3[17]), .sel(shft[3]), 
      .out(z4[17]));
   mux2X1_r__0_433 genblk1_11_m8 (.in0(z3[24]), .in1(z3[16]), .sel(shft[3]), 
      .out(z4[16]));
   mux2X1_r__0_435 genblk1_12_m8 (.in0(z3[23]), .in1(z3[15]), .sel(shft[3]), 
      .out(z4[15]));
   mux2X1_r__0_437 genblk1_13_m8 (.in0(z3[22]), .in1(z3[14]), .sel(shft[3]), 
      .out(z4[14]));
   mux2X1_r__0_439 genblk1_14_m8 (.in0(z3[21]), .in1(z3[13]), .sel(shft[3]), 
      .out(z4[13]));
   mux2X1_r__0_441 genblk1_15_m8 (.in0(z3[20]), .in1(z3[12]), .sel(shft[3]), 
      .out(z4[12]));
   mux2X1_r__0_443 genblk1_16_m8 (.in0(z3[19]), .in1(z3[11]), .sel(shft[3]), 
      .out(z4[11]));
   mux2X1_r__0_445 genblk1_17_m8 (.in0(z3[18]), .in1(z3[10]), .sel(shft[3]), 
      .out(z4[10]));
   mux2X1_r__0_447 genblk1_18_m8 (.in0(z3[17]), .in1(z3[9]), .sel(shft[3]), 
      .out(z4[9]));
   mux2X1_r__0_449 genblk1_19_m8 (.in0(z3[16]), .in1(z3[8]), .sel(shft[3]), 
      .out(z4[8]));
   mux2X1_r__0_451 genblk1_20_m8 (.in0(z3[15]), .in1(z3[7]), .sel(shft[3]), 
      .out(z4[7]));
   mux2X1_r__0_453 genblk1_21_m8 (.in0(z3[14]), .in1(z3[6]), .sel(shft[3]), 
      .out(z4[6]));
   mux2X1_r__0_455 genblk1_22_m8 (.in0(z3[13]), .in1(z3[5]), .sel(shft[3]), 
      .out(z4[5]));
   mux2X1_r__0_457 genblk1_23_m8 (.in0(z3[12]), .in1(z3[4]), .sel(shft[3]), 
      .out(z4[4]));
   mux2X1_r__0_459 genblk1_24_m8 (.in0(z3[11]), .in1(z3[3]), .sel(shft[3]), 
      .out(z4[3]));
   mux2X1_r__0_461 genblk1_25_m8 (.in0(z3[10]), .in1(z3[2]), .sel(shft[3]), 
      .out(z4[2]));
   mux2X1_r__0_463 genblk1_26_m8 (.in0(z3[9]), .in1(z3[1]), .sel(shft[3]), 
      .out(z4[1]));
   mux2X1_r__0_465 genblk1_27_m8 (.in0(z3[8]), .in1(z3[0]), .sel(shft[3]), 
      .out(z4[0]));
   mux2X1_r__0_467 genblk1_0_m5 (.in0(), .in1(z2[27]), .sel(shft[2]), .out(
      z3[27]));
   mux2X1_r__0_469 genblk1_1_m5 (.in0(), .in1(z2[26]), .sel(shft[2]), .out(
      z3[26]));
   mux2X1_r__0_471 genblk1_2_m5 (.in0(), .in1(z2[25]), .sel(shft[2]), .out(
      z3[25]));
   mux2X1_r__0_473 genblk1_3_m5 (.in0(), .in1(z2[24]), .sel(shft[2]), .out(
      z3[24]));
   mux2X1_r__0_475 genblk1_4_m6 (.in0(z2[27]), .in1(z2[23]), .sel(shft[2]), 
      .out(z3[23]));
   mux2X1_r__0_477 genblk1_5_m6 (.in0(z2[26]), .in1(z2[22]), .sel(shft[2]), 
      .out(z3[22]));
   mux2X1_r__0_479 genblk1_6_m6 (.in0(z2[25]), .in1(z2[21]), .sel(shft[2]), 
      .out(z3[21]));
   mux2X1_r__0_481 genblk1_7_m6 (.in0(z2[24]), .in1(z2[20]), .sel(shft[2]), 
      .out(z3[20]));
   mux2X1_r__0_483 genblk1_8_m6 (.in0(z2[23]), .in1(z2[19]), .sel(shft[2]), 
      .out(z3[19]));
   mux2X1_r__0_485 genblk1_9_m6 (.in0(z2[22]), .in1(z2[18]), .sel(shft[2]), 
      .out(z3[18]));
   mux2X1_r__0_487 genblk1_10_m6 (.in0(z2[21]), .in1(z2[17]), .sel(shft[2]), 
      .out(z3[17]));
   mux2X1_r__0_489 genblk1_11_m6 (.in0(z2[20]), .in1(z2[16]), .sel(shft[2]), 
      .out(z3[16]));
   mux2X1_r__0_491 genblk1_12_m6 (.in0(z2[19]), .in1(z2[15]), .sel(shft[2]), 
      .out(z3[15]));
   mux2X1_r__0_493 genblk1_13_m6 (.in0(z2[18]), .in1(z2[14]), .sel(shft[2]), 
      .out(z3[14]));
   mux2X1_r__0_495 genblk1_14_m6 (.in0(z2[17]), .in1(z2[13]), .sel(shft[2]), 
      .out(z3[13]));
   mux2X1_r__0_497 genblk1_15_m6 (.in0(z2[16]), .in1(z2[12]), .sel(shft[2]), 
      .out(z3[12]));
   mux2X1_r__0_499 genblk1_16_m6 (.in0(z2[15]), .in1(z2[11]), .sel(shft[2]), 
      .out(z3[11]));
   mux2X1_r__0_501 genblk1_17_m6 (.in0(z2[14]), .in1(z2[10]), .sel(shft[2]), 
      .out(z3[10]));
   mux2X1_r__0_503 genblk1_18_m6 (.in0(z2[13]), .in1(z2[9]), .sel(shft[2]), 
      .out(z3[9]));
   mux2X1_r__0_505 genblk1_19_m6 (.in0(z2[12]), .in1(z2[8]), .sel(shft[2]), 
      .out(z3[8]));
   mux2X1_r__0_507 genblk1_20_m6 (.in0(z2[11]), .in1(z2[7]), .sel(shft[2]), 
      .out(z3[7]));
   mux2X1_r__0_509 genblk1_21_m6 (.in0(z2[10]), .in1(z2[6]), .sel(shft[2]), 
      .out(z3[6]));
   mux2X1_r__0_511 genblk1_22_m6 (.in0(z2[9]), .in1(z2[5]), .sel(shft[2]), 
      .out(z3[5]));
   mux2X1_r__0_513 genblk1_23_m6 (.in0(z2[8]), .in1(z2[4]), .sel(shft[2]), 
      .out(z3[4]));
   mux2X1_r__0_515 genblk1_24_m6 (.in0(z2[7]), .in1(z2[3]), .sel(shft[2]), 
      .out(z3[3]));
   mux2X1_r__0_517 genblk1_25_m6 (.in0(z2[6]), .in1(z2[2]), .sel(shft[2]), 
      .out(z3[2]));
   mux2X1_r__0_519 genblk1_26_m6 (.in0(z2[5]), .in1(z2[1]), .sel(shft[2]), 
      .out(z3[1]));
   mux2X1_r__0_521 genblk1_27_m6 (.in0(z2[4]), .in1(), .sel(shft[2]), .out(z3[0]));
   mux2X1_r__0_523 genblk1_0_m3 (.in0(), .in1(z1[27]), .sel(shft[1]), .out(
      z2[27]));
   mux2X1_r__0_525 genblk1_1_m3 (.in0(), .in1(z1[26]), .sel(shft[1]), .out(
      z2[26]));
   mux2X1_r__0_527 genblk1_2_m4 (.in0(z1[27]), .in1(z1[25]), .sel(shft[1]), 
      .out(z2[25]));
   mux2X1_r__0_529 genblk1_3_m4 (.in0(z1[26]), .in1(z1[24]), .sel(shft[1]), 
      .out(z2[24]));
   mux2X1_r__0_531 genblk1_4_m4 (.in0(z1[25]), .in1(z1[23]), .sel(shft[1]), 
      .out(z2[23]));
   mux2X1_r__0_533 genblk1_5_m4 (.in0(z1[24]), .in1(z1[22]), .sel(shft[1]), 
      .out(z2[22]));
   mux2X1_r__0_535 genblk1_6_m4 (.in0(z1[23]), .in1(z1[21]), .sel(shft[1]), 
      .out(z2[21]));
   mux2X1_r__0_537 genblk1_7_m4 (.in0(z1[22]), .in1(z1[20]), .sel(shft[1]), 
      .out(z2[20]));
   mux2X1_r__0_539 genblk1_8_m4 (.in0(z1[21]), .in1(z1[19]), .sel(shft[1]), 
      .out(z2[19]));
   mux2X1_r__0_541 genblk1_9_m4 (.in0(z1[20]), .in1(z1[18]), .sel(shft[1]), 
      .out(z2[18]));
   mux2X1_r__0_543 genblk1_10_m4 (.in0(z1[19]), .in1(z1[17]), .sel(shft[1]), 
      .out(z2[17]));
   mux2X1_r__0_545 genblk1_11_m4 (.in0(z1[18]), .in1(z1[16]), .sel(shft[1]), 
      .out(z2[16]));
   mux2X1_r__0_547 genblk1_12_m4 (.in0(z1[17]), .in1(z1[15]), .sel(shft[1]), 
      .out(z2[15]));
   mux2X1_r__0_549 genblk1_13_m4 (.in0(z1[16]), .in1(z1[14]), .sel(shft[1]), 
      .out(z2[14]));
   mux2X1_r__0_551 genblk1_14_m4 (.in0(z1[15]), .in1(z1[13]), .sel(shft[1]), 
      .out(z2[13]));
   mux2X1_r__0_553 genblk1_15_m4 (.in0(z1[14]), .in1(z1[12]), .sel(shft[1]), 
      .out(z2[12]));
   mux2X1_r__0_555 genblk1_16_m4 (.in0(z1[13]), .in1(z1[11]), .sel(shft[1]), 
      .out(z2[11]));
   mux2X1_r__0_557 genblk1_17_m4 (.in0(z1[12]), .in1(z1[10]), .sel(shft[1]), 
      .out(z2[10]));
   mux2X1_r__0_559 genblk1_18_m4 (.in0(z1[11]), .in1(z1[9]), .sel(shft[1]), 
      .out(z2[9]));
   mux2X1_r__0_561 genblk1_19_m4 (.in0(z1[10]), .in1(z1[8]), .sel(shft[1]), 
      .out(z2[8]));
   mux2X1_r__0_563 genblk1_20_m4 (.in0(z1[9]), .in1(z1[7]), .sel(shft[1]), 
      .out(z2[7]));
   mux2X1_r__0_565 genblk1_21_m4 (.in0(z1[8]), .in1(z1[6]), .sel(shft[1]), 
      .out(z2[6]));
   mux2X1_r__0_567 genblk1_22_m4 (.in0(z1[7]), .in1(z1[5]), .sel(shft[1]), 
      .out(z2[5]));
   mux2X1_r__0_569 genblk1_23_m4 (.in0(z1[6]), .in1(z1[4]), .sel(shft[1]), 
      .out(z2[4]));
   mux2X1_r__0_571 genblk1_24_m4 (.in0(z1[5]), .in1(z1[3]), .sel(shft[1]), 
      .out(z2[3]));
   mux2X1_r__0_573 genblk1_25_m4 (.in0(z1[4]), .in1(), .sel(shft[1]), .out(z2[2]));
   mux2X1_r__0_575 genblk1_26_m4 (.in0(z1[3]), .in1(), .sel(shft[1]), .out(z2[1]));
   mux2X1_r__0_579 genblk1_0_m1 (.in0(), .in1(in[27]), .sel(shft[0]), .out(
      z1[27]));
   mux2X1_r__0_581 genblk1_1_m2 (.in0(in[27]), .in1(in[26]), .sel(shft[0]), 
      .out(z1[26]));
   mux2X1_r__0_583 genblk1_2_m2 (.in0(in[26]), .in1(in[25]), .sel(shft[0]), 
      .out(z1[25]));
   mux2X1_r__0_585 genblk1_3_m2 (.in0(in[25]), .in1(in[24]), .sel(shft[0]), 
      .out(z1[24]));
   mux2X1_r__0_587 genblk1_4_m2 (.in0(in[24]), .in1(in[23]), .sel(shft[0]), 
      .out(z1[23]));
   mux2X1_r__0_589 genblk1_5_m2 (.in0(in[23]), .in1(in[22]), .sel(shft[0]), 
      .out(z1[22]));
   mux2X1_r__0_591 genblk1_6_m2 (.in0(in[22]), .in1(in[21]), .sel(shft[0]), 
      .out(z1[21]));
   mux2X1_r__0_593 genblk1_7_m2 (.in0(in[21]), .in1(in[20]), .sel(shft[0]), 
      .out(z1[20]));
   mux2X1_r__0_595 genblk1_8_m2 (.in0(in[20]), .in1(in[19]), .sel(shft[0]), 
      .out(z1[19]));
   mux2X1_r__0_597 genblk1_9_m2 (.in0(in[19]), .in1(in[18]), .sel(shft[0]), 
      .out(z1[18]));
   mux2X1_r__0_599 genblk1_10_m2 (.in0(in[18]), .in1(in[17]), .sel(shft[0]), 
      .out(z1[17]));
   mux2X1_r__0_601 genblk1_11_m2 (.in0(in[17]), .in1(in[16]), .sel(shft[0]), 
      .out(z1[16]));
   mux2X1_r__0_603 genblk1_12_m2 (.in0(in[16]), .in1(in[15]), .sel(shft[0]), 
      .out(z1[15]));
   mux2X1_r__0_605 genblk1_13_m2 (.in0(in[15]), .in1(in[14]), .sel(shft[0]), 
      .out(z1[14]));
   mux2X1_r__0_607 genblk1_14_m2 (.in0(in[14]), .in1(in[13]), .sel(shft[0]), 
      .out(z1[13]));
   mux2X1_r__0_609 genblk1_15_m2 (.in0(in[13]), .in1(in[12]), .sel(shft[0]), 
      .out(z1[12]));
   mux2X1_r__0_611 genblk1_16_m2 (.in0(in[12]), .in1(in[11]), .sel(shft[0]), 
      .out(z1[11]));
   mux2X1_r__0_613 genblk1_17_m2 (.in0(in[11]), .in1(in[10]), .sel(shft[0]), 
      .out(z1[10]));
   mux2X1_r__0_615 genblk1_18_m2 (.in0(in[10]), .in1(in[9]), .sel(shft[0]), 
      .out(z1[9]));
   mux2X1_r__0_617 genblk1_19_m2 (.in0(in[9]), .in1(in[8]), .sel(shft[0]), 
      .out(z1[8]));
   mux2X1_r__0_619 genblk1_20_m2 (.in0(in[8]), .in1(in[7]), .sel(shft[0]), 
      .out(z1[7]));
   mux2X1_r__0_621 genblk1_21_m2 (.in0(in[7]), .in1(in[6]), .sel(shft[0]), 
      .out(z1[6]));
   mux2X1_r__0_623 genblk1_22_m2 (.in0(in[6]), .in1(in[5]), .sel(shft[0]), 
      .out(z1[5]));
   mux2X1_r__0_625 genblk1_23_m2 (.in0(in[5]), .in1(in[4]), .sel(shft[0]), 
      .out(z1[4]));
   mux2X1_r__0_627 genblk1_24_m2 (.in0(in[4]), .in1(), .sel(shft[0]), .out(z1[3]));
endmodule

module n_normal(A, B, edata, SA, SB, Comp, Enor, MA, MB);
   input [36:0]A;
   input [36:0]B;
   input [1:0]edata;
   output SA;
   output SB;
   output Comp;
   output [7:0]Enor;
   output [27:0]MA;
   output [27:0]MB;

   wire [4:0]Dexp;
   wire [27:0]MShift;

   comp_exp com (.A({uc_0, A[35], A[34], A[33], A[32], A[31], A[30], A[29], 
      A[28], A[27], A[26], A[25], A[24], A[23], A[22], A[21], A[20], A[19], 
      A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], 
      A[7], A[6], A[5], A[4], uc_1, uc_2, uc_3, uc_4}), .B({uc_5, B[35], B[34], 
      B[33], B[32], B[31], B[30], B[29], B[28], B[27], B[26], B[25], B[24], 
      B[23], B[22], B[21], B[20], B[19], B[18], B[17], B[16], B[15], B[14], 
      B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], B[5], B[4], uc_6, uc_7, 
      uc_8, uc_9}), .edata(edata), .SA(), .SB(), .Comp(Comp), .Enor(Enor), 
      .MMax({MA[27], MA[26], MA[25], MA[24], MA[23], MA[22], MA[21], MA[20], 
      MA[19], MA[18], MA[17], MA[16], MA[15], MA[14], MA[13], MA[12], MA[11], 
      MA[10], MA[9], MA[8], MA[7], MA[6], MA[5], MA[4], uc_10, uc_11, uc_12, 
      uc_13}), .MShift({MShift[27], MShift[26], MShift[25], MShift[24], 
      MShift[23], MShift[22], MShift[21], MShift[20], MShift[19], MShift[18], 
      MShift[17], MShift[16], MShift[15], MShift[14], MShift[13], MShift[12], 
      MShift[11], MShift[10], MShift[9], MShift[8], MShift[7], MShift[6], 
      MShift[5], MShift[4], uc_14, uc_15, uc_16, uc_17}), .Dexp(Dexp));
   n_shift_norm sh (.shft(Dexp), .in({MShift[27], MShift[26], MShift[25], 
      MShift[24], MShift[23], MShift[22], MShift[21], MShift[20], MShift[19], 
      MShift[18], MShift[17], MShift[16], MShift[15], MShift[14], MShift[13], 
      MShift[12], MShift[11], MShift[10], MShift[9], MShift[8], MShift[7], 
      MShift[6], MShift[5], MShift[4], uc_18, uc_19, uc_20, uc_21}), .out(MB));
endmodule

module mux_adder(SAsub, SBsub, SComp, Esub, MAsub, MBsub, SAnor, SBnor, NComp, 
      Enor, MAnor, MBnor, edata, SA, SB, C, Eout, MAout, MBout);
   input SAsub;
   input SBsub;
   input SComp;
   input [7:0]Esub;
   input [27:0]MAsub;
   input [27:0]MBsub;
   input SAnor;
   input SBnor;
   input NComp;
   input [7:0]Enor;
   input [27:0]MAnor;
   input [27:0]MBnor;
   input [1:0]edata;
   output SA;
   output SB;
   output C;
   output [7:0]Eout;
   output [27:0]MAout;
   output [27:0]MBout;

   wire n_0_0;

   OR2_X1 i_0_0 (.A1(edata[1]), .A2(edata[0]), .ZN(n_0_0));
   MUX2_X1 i_0_1 (.A(SComp), .B(NComp), .S(n_0_0), .Z(C));
   MUX2_X1 i_0_2 (.A(Esub[0]), .B(Enor[0]), .S(n_0_0), .Z(Eout[0]));
   MUX2_X1 i_0_3 (.A(Esub[1]), .B(Enor[1]), .S(n_0_0), .Z(Eout[1]));
   MUX2_X1 i_0_4 (.A(Esub[2]), .B(Enor[2]), .S(n_0_0), .Z(Eout[2]));
   MUX2_X1 i_0_5 (.A(Esub[3]), .B(Enor[3]), .S(n_0_0), .Z(Eout[3]));
   MUX2_X1 i_0_6 (.A(Esub[4]), .B(Enor[4]), .S(n_0_0), .Z(Eout[4]));
   MUX2_X1 i_0_7 (.A(Esub[5]), .B(Enor[5]), .S(n_0_0), .Z(Eout[5]));
   MUX2_X1 i_0_8 (.A(Esub[6]), .B(Enor[6]), .S(n_0_0), .Z(Eout[6]));
   MUX2_X1 i_0_9 (.A(Esub[7]), .B(Enor[7]), .S(n_0_0), .Z(Eout[7]));
   MUX2_X1 i_0_10 (.A(MAsub[4]), .B(MAnor[4]), .S(n_0_0), .Z(MAout[4]));
   MUX2_X1 i_0_11 (.A(MAsub[5]), .B(MAnor[5]), .S(n_0_0), .Z(MAout[5]));
   MUX2_X1 i_0_12 (.A(MAsub[6]), .B(MAnor[6]), .S(n_0_0), .Z(MAout[6]));
   MUX2_X1 i_0_13 (.A(MAsub[7]), .B(MAnor[7]), .S(n_0_0), .Z(MAout[7]));
   MUX2_X1 i_0_14 (.A(MAsub[8]), .B(MAnor[8]), .S(n_0_0), .Z(MAout[8]));
   MUX2_X1 i_0_15 (.A(MAsub[9]), .B(MAnor[9]), .S(n_0_0), .Z(MAout[9]));
   MUX2_X1 i_0_16 (.A(MAsub[10]), .B(MAnor[10]), .S(n_0_0), .Z(MAout[10]));
   MUX2_X1 i_0_17 (.A(MAsub[11]), .B(MAnor[11]), .S(n_0_0), .Z(MAout[11]));
   MUX2_X1 i_0_18 (.A(MAsub[12]), .B(MAnor[12]), .S(n_0_0), .Z(MAout[12]));
   MUX2_X1 i_0_19 (.A(MAsub[13]), .B(MAnor[13]), .S(n_0_0), .Z(MAout[13]));
   MUX2_X1 i_0_20 (.A(MAsub[14]), .B(MAnor[14]), .S(n_0_0), .Z(MAout[14]));
   MUX2_X1 i_0_21 (.A(MAsub[15]), .B(MAnor[15]), .S(n_0_0), .Z(MAout[15]));
   MUX2_X1 i_0_22 (.A(MAsub[16]), .B(MAnor[16]), .S(n_0_0), .Z(MAout[16]));
   MUX2_X1 i_0_23 (.A(MAsub[17]), .B(MAnor[17]), .S(n_0_0), .Z(MAout[17]));
   MUX2_X1 i_0_24 (.A(MAsub[18]), .B(MAnor[18]), .S(n_0_0), .Z(MAout[18]));
   MUX2_X1 i_0_25 (.A(MAsub[19]), .B(MAnor[19]), .S(n_0_0), .Z(MAout[19]));
   MUX2_X1 i_0_26 (.A(MAsub[20]), .B(MAnor[20]), .S(n_0_0), .Z(MAout[20]));
   MUX2_X1 i_0_27 (.A(MAsub[21]), .B(MAnor[21]), .S(n_0_0), .Z(MAout[21]));
   MUX2_X1 i_0_28 (.A(MAsub[22]), .B(MAnor[22]), .S(n_0_0), .Z(MAout[22]));
   MUX2_X1 i_0_29 (.A(MAsub[23]), .B(MAnor[23]), .S(n_0_0), .Z(MAout[23]));
   MUX2_X1 i_0_30 (.A(MAsub[24]), .B(MAnor[24]), .S(n_0_0), .Z(MAout[24]));
   MUX2_X1 i_0_31 (.A(MAsub[25]), .B(MAnor[25]), .S(n_0_0), .Z(MAout[25]));
   MUX2_X1 i_0_32 (.A(MAsub[26]), .B(MAnor[26]), .S(n_0_0), .Z(MAout[26]));
   MUX2_X1 i_0_33 (.A(MAsub[27]), .B(MAnor[27]), .S(n_0_0), .Z(MAout[27]));
   AND2_X1 i_0_34 (.A1(n_0_0), .A2(MBnor[0]), .ZN(MBout[0]));
   AND2_X1 i_0_35 (.A1(n_0_0), .A2(MBnor[1]), .ZN(MBout[1]));
   AND2_X1 i_0_36 (.A1(n_0_0), .A2(MBnor[2]), .ZN(MBout[2]));
   AND2_X1 i_0_37 (.A1(n_0_0), .A2(MBnor[3]), .ZN(MBout[3]));
   MUX2_X1 i_0_38 (.A(MBsub[4]), .B(MBnor[4]), .S(n_0_0), .Z(MBout[4]));
   MUX2_X1 i_0_39 (.A(MBsub[5]), .B(MBnor[5]), .S(n_0_0), .Z(MBout[5]));
   MUX2_X1 i_0_40 (.A(MBsub[6]), .B(MBnor[6]), .S(n_0_0), .Z(MBout[6]));
   MUX2_X1 i_0_41 (.A(MBsub[7]), .B(MBnor[7]), .S(n_0_0), .Z(MBout[7]));
   MUX2_X1 i_0_42 (.A(MBsub[8]), .B(MBnor[8]), .S(n_0_0), .Z(MBout[8]));
   MUX2_X1 i_0_43 (.A(MBsub[9]), .B(MBnor[9]), .S(n_0_0), .Z(MBout[9]));
   MUX2_X1 i_0_44 (.A(MBsub[10]), .B(MBnor[10]), .S(n_0_0), .Z(MBout[10]));
   MUX2_X1 i_0_45 (.A(MBsub[11]), .B(MBnor[11]), .S(n_0_0), .Z(MBout[11]));
   MUX2_X1 i_0_46 (.A(MBsub[12]), .B(MBnor[12]), .S(n_0_0), .Z(MBout[12]));
   MUX2_X1 i_0_47 (.A(MBsub[13]), .B(MBnor[13]), .S(n_0_0), .Z(MBout[13]));
   MUX2_X1 i_0_48 (.A(MBsub[14]), .B(MBnor[14]), .S(n_0_0), .Z(MBout[14]));
   MUX2_X1 i_0_49 (.A(MBsub[15]), .B(MBnor[15]), .S(n_0_0), .Z(MBout[15]));
   MUX2_X1 i_0_50 (.A(MBsub[16]), .B(MBnor[16]), .S(n_0_0), .Z(MBout[16]));
   MUX2_X1 i_0_51 (.A(MBsub[17]), .B(MBnor[17]), .S(n_0_0), .Z(MBout[17]));
   MUX2_X1 i_0_52 (.A(MBsub[18]), .B(MBnor[18]), .S(n_0_0), .Z(MBout[18]));
   MUX2_X1 i_0_53 (.A(MBsub[19]), .B(MBnor[19]), .S(n_0_0), .Z(MBout[19]));
   MUX2_X1 i_0_54 (.A(MBsub[20]), .B(MBnor[20]), .S(n_0_0), .Z(MBout[20]));
   MUX2_X1 i_0_55 (.A(MBsub[21]), .B(MBnor[21]), .S(n_0_0), .Z(MBout[21]));
   MUX2_X1 i_0_56 (.A(MBsub[22]), .B(MBnor[22]), .S(n_0_0), .Z(MBout[22]));
   MUX2_X1 i_0_57 (.A(MBsub[23]), .B(MBnor[23]), .S(n_0_0), .Z(MBout[23]));
   MUX2_X1 i_0_58 (.A(MBsub[24]), .B(MBnor[24]), .S(n_0_0), .Z(MBout[24]));
   MUX2_X1 i_0_59 (.A(MBsub[25]), .B(MBnor[25]), .S(n_0_0), .Z(MBout[25]));
   MUX2_X1 i_0_60 (.A(MBsub[26]), .B(MBnor[26]), .S(n_0_0), .Z(MBout[26]));
   MUX2_X1 i_0_61 (.A(MBsub[27]), .B(MBnor[27]), .S(n_0_0), .Z(MBout[27]));
endmodule

module signout(SA, SB, Comp, A, B, A_S, Aa, Bb, AS, SO);
   input SA;
   input SB;
   input Comp;
   input [27:0]A;
   input [27:0]B;
   input A_S;
   output [27:0]Aa;
   output [27:0]Bb;
   output AS;
   output SO;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_3), .B2(Comp), .ZN(SO));
   NAND2_X1 i_0_1 (.A1(SA), .A2(Comp), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(B[0]), .A2(n_0_1), .ZN(Bb[0]));
   AND2_X1 i_0_3 (.A1(B[1]), .A2(n_0_1), .ZN(Bb[1]));
   AND2_X1 i_0_4 (.A1(B[2]), .A2(n_0_1), .ZN(Bb[2]));
   AND2_X1 i_0_5 (.A1(B[3]), .A2(n_0_1), .ZN(Bb[3]));
   MUX2_X1 i_0_6 (.A(A[4]), .B(B[4]), .S(n_0_1), .Z(Bb[4]));
   MUX2_X1 i_0_7 (.A(A[5]), .B(B[5]), .S(n_0_1), .Z(Bb[5]));
   MUX2_X1 i_0_8 (.A(A[6]), .B(B[6]), .S(n_0_1), .Z(Bb[6]));
   MUX2_X1 i_0_9 (.A(A[7]), .B(B[7]), .S(n_0_1), .Z(Bb[7]));
   MUX2_X1 i_0_10 (.A(A[8]), .B(B[8]), .S(n_0_1), .Z(Bb[8]));
   MUX2_X1 i_0_11 (.A(A[9]), .B(B[9]), .S(n_0_1), .Z(Bb[9]));
   MUX2_X1 i_0_12 (.A(A[10]), .B(B[10]), .S(n_0_1), .Z(Bb[10]));
   MUX2_X1 i_0_13 (.A(A[11]), .B(B[11]), .S(n_0_1), .Z(Bb[11]));
   MUX2_X1 i_0_14 (.A(A[12]), .B(B[12]), .S(n_0_1), .Z(Bb[12]));
   MUX2_X1 i_0_15 (.A(A[13]), .B(B[13]), .S(n_0_1), .Z(Bb[13]));
   MUX2_X1 i_0_16 (.A(A[14]), .B(B[14]), .S(n_0_1), .Z(Bb[14]));
   MUX2_X1 i_0_17 (.A(A[15]), .B(B[15]), .S(n_0_1), .Z(Bb[15]));
   MUX2_X1 i_0_18 (.A(A[16]), .B(B[16]), .S(n_0_1), .Z(Bb[16]));
   MUX2_X1 i_0_19 (.A(A[17]), .B(B[17]), .S(n_0_1), .Z(Bb[17]));
   MUX2_X1 i_0_20 (.A(A[18]), .B(B[18]), .S(n_0_1), .Z(Bb[18]));
   MUX2_X1 i_0_21 (.A(A[19]), .B(B[19]), .S(n_0_1), .Z(Bb[19]));
   MUX2_X1 i_0_22 (.A(A[20]), .B(B[20]), .S(n_0_1), .Z(Bb[20]));
   MUX2_X1 i_0_23 (.A(A[21]), .B(B[21]), .S(n_0_1), .Z(Bb[21]));
   MUX2_X1 i_0_24 (.A(A[22]), .B(B[22]), .S(n_0_1), .Z(Bb[22]));
   MUX2_X1 i_0_25 (.A(A[23]), .B(B[23]), .S(n_0_1), .Z(Bb[23]));
   MUX2_X1 i_0_26 (.A(A[24]), .B(B[24]), .S(n_0_1), .Z(Bb[24]));
   MUX2_X1 i_0_27 (.A(A[25]), .B(B[25]), .S(n_0_1), .Z(Bb[25]));
   MUX2_X1 i_0_28 (.A(A[26]), .B(B[26]), .S(n_0_1), .Z(Bb[26]));
   MUX2_X1 i_0_29 (.A(A[27]), .B(B[27]), .S(n_0_1), .Z(Bb[27]));
   AND2_X1 i_0_30 (.A1(n_0_4), .A2(B[0]), .ZN(Aa[0]));
   AND2_X1 i_0_31 (.A1(n_0_4), .A2(B[1]), .ZN(Aa[1]));
   AND2_X1 i_0_32 (.A1(n_0_4), .A2(B[2]), .ZN(Aa[2]));
   AND2_X1 i_0_33 (.A1(n_0_4), .A2(B[3]), .ZN(Aa[3]));
   MUX2_X1 i_0_34 (.A(B[4]), .B(A[4]), .S(n_0_1), .Z(Aa[4]));
   MUX2_X1 i_0_35 (.A(B[5]), .B(A[5]), .S(n_0_1), .Z(Aa[5]));
   MUX2_X1 i_0_36 (.A(B[6]), .B(A[6]), .S(n_0_1), .Z(Aa[6]));
   MUX2_X1 i_0_37 (.A(B[7]), .B(A[7]), .S(n_0_1), .Z(Aa[7]));
   MUX2_X1 i_0_38 (.A(B[8]), .B(A[8]), .S(n_0_1), .Z(Aa[8]));
   MUX2_X1 i_0_39 (.A(B[9]), .B(A[9]), .S(n_0_1), .Z(Aa[9]));
   MUX2_X1 i_0_40 (.A(B[10]), .B(A[10]), .S(n_0_1), .Z(Aa[10]));
   MUX2_X1 i_0_41 (.A(B[11]), .B(A[11]), .S(n_0_1), .Z(Aa[11]));
   MUX2_X1 i_0_42 (.A(B[12]), .B(A[12]), .S(n_0_1), .Z(Aa[12]));
   MUX2_X1 i_0_43 (.A(B[13]), .B(A[13]), .S(n_0_1), .Z(Aa[13]));
   MUX2_X1 i_0_44 (.A(B[14]), .B(A[14]), .S(n_0_1), .Z(Aa[14]));
   MUX2_X1 i_0_45 (.A(B[15]), .B(A[15]), .S(n_0_1), .Z(Aa[15]));
   MUX2_X1 i_0_46 (.A(B[16]), .B(A[16]), .S(n_0_1), .Z(Aa[16]));
   MUX2_X1 i_0_47 (.A(B[17]), .B(A[17]), .S(n_0_1), .Z(Aa[17]));
   MUX2_X1 i_0_48 (.A(B[18]), .B(A[18]), .S(n_0_1), .Z(Aa[18]));
   MUX2_X1 i_0_49 (.A(B[19]), .B(A[19]), .S(n_0_1), .Z(Aa[19]));
   MUX2_X1 i_0_50 (.A(B[20]), .B(A[20]), .S(n_0_1), .Z(Aa[20]));
   MUX2_X1 i_0_51 (.A(B[21]), .B(A[21]), .S(n_0_1), .Z(Aa[21]));
   MUX2_X1 i_0_52 (.A(B[22]), .B(A[22]), .S(n_0_1), .Z(Aa[22]));
   MUX2_X1 i_0_53 (.A(B[23]), .B(A[23]), .S(n_0_1), .Z(Aa[23]));
   MUX2_X1 i_0_54 (.A(B[24]), .B(A[24]), .S(n_0_1), .Z(Aa[24]));
   MUX2_X1 i_0_55 (.A(B[25]), .B(A[25]), .S(n_0_1), .Z(Aa[25]));
   MUX2_X1 i_0_56 (.A(B[26]), .B(A[26]), .S(n_0_1), .Z(Aa[26]));
   MUX2_X1 i_0_57 (.A(B[27]), .B(A[27]), .S(n_0_1), .Z(Aa[27]));
   XNOR2_X1 i_0_58 (.A(Comp), .B(n_0_2), .ZN(n_0_1));
   XNOR2_X1 i_0_59 (.A(SA), .B(n_0_3), .ZN(AS));
   NAND2_X1 i_0_60 (.A1(n_0_3), .A2(SA), .ZN(n_0_2));
   XNOR2_X1 i_0_61 (.A(A_S), .B(SB), .ZN(n_0_3));
   INV_X1 i_0_62 (.A(n_0_1), .ZN(n_0_4));
endmodule

module datapath__0_54(add1_i, p_0, add2_i);
   input [27:0]add1_i;
   output [28:0]p_0;
   input [27:0]add2_i;

   INV_X1 i_0 (.A(add1_i[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(add2_i[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(add2_i[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(add1_i[1]), .B(add2_i[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(add1_i[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(add2_i[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(add1_i[2]), .B(add2_i[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(add2_i[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(add1_i[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(add1_i[3]), .B(add2_i[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(add1_i[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(add2_i[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(add1_i[4]), .B(add2_i[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(add2_i[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(add1_i[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(add1_i[5]), .B(add2_i[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(add1_i[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(add2_i[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(add1_i[6]), .B(add2_i[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(add2_i[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(add1_i[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(add1_i[7]), .B(add2_i[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(add1_i[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(add2_i[7]), .ZN(n_23));
   INV_X1 i_32 (.A(add1_i[8]), .ZN(n_24));
   OR2_X1 i_33 (.A1(n_24), .A2(add2_i[8]), .ZN(n_25));
   NAND2_X1 i_34 (.A1(n_24), .A2(add2_i[8]), .ZN(n_26));
   NAND2_X1 i_35 (.A1(n_25), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_36 (.A(n_23), .B(n_27), .ZN(p_0[8]));
   INV_X1 i_37 (.A(n_25), .ZN(n_28));
   AOI21_X1 i_38 (.A(n_28), .B1(n_23), .B2(n_26), .ZN(n_29));
   XNOR2_X1 i_39 (.A(add1_i[9]), .B(add2_i[9]), .ZN(n_30));
   XNOR2_X1 i_40 (.A(n_29), .B(n_30), .ZN(p_0[9]));
   INV_X1 i_41 (.A(add1_i[9]), .ZN(n_31));
   AOI22_X1 i_42 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(add2_i[9]), .ZN(n_32));
   XOR2_X1 i_43 (.A(add1_i[10]), .B(add2_i[10]), .Z(n_33));
   XNOR2_X1 i_44 (.A(n_32), .B(n_33), .ZN(p_0[10]));
   INV_X1 i_45 (.A(add2_i[10]), .ZN(n_34));
   OAI22_X1 i_46 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(add1_i[10]), .ZN(n_35));
   XNOR2_X1 i_47 (.A(add1_i[11]), .B(add2_i[11]), .ZN(n_36));
   XNOR2_X1 i_48 (.A(n_35), .B(n_36), .ZN(p_0[11]));
   INV_X1 i_49 (.A(add1_i[11]), .ZN(n_37));
   AOI22_X1 i_50 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(add2_i[11]), .ZN(n_38));
   XOR2_X1 i_51 (.A(add1_i[12]), .B(add2_i[12]), .Z(n_39));
   XNOR2_X1 i_52 (.A(n_38), .B(n_39), .ZN(p_0[12]));
   INV_X1 i_53 (.A(add2_i[12]), .ZN(n_40));
   OAI22_X1 i_54 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(add1_i[12]), .ZN(n_41));
   XNOR2_X1 i_55 (.A(add1_i[13]), .B(add2_i[13]), .ZN(n_42));
   XNOR2_X1 i_56 (.A(n_41), .B(n_42), .ZN(p_0[13]));
   INV_X1 i_57 (.A(add1_i[13]), .ZN(n_43));
   AOI22_X1 i_58 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(add2_i[13]), .ZN(n_44));
   XOR2_X1 i_59 (.A(add1_i[14]), .B(add2_i[14]), .Z(n_45));
   XNOR2_X1 i_60 (.A(n_44), .B(n_45), .ZN(p_0[14]));
   INV_X1 i_61 (.A(add2_i[14]), .ZN(n_46));
   OAI22_X1 i_62 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(add1_i[14]), .ZN(n_47));
   XNOR2_X1 i_63 (.A(add1_i[15]), .B(add2_i[15]), .ZN(n_48));
   XNOR2_X1 i_64 (.A(n_47), .B(n_48), .ZN(p_0[15]));
   INV_X1 i_65 (.A(add1_i[15]), .ZN(n_49));
   AOI22_X1 i_66 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(add2_i[15]), .ZN(n_50));
   XOR2_X1 i_67 (.A(add1_i[16]), .B(add2_i[16]), .Z(n_51));
   XNOR2_X1 i_68 (.A(n_50), .B(n_51), .ZN(p_0[16]));
   INV_X1 i_69 (.A(add2_i[16]), .ZN(n_52));
   OAI22_X1 i_70 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(add1_i[16]), .ZN(n_53));
   XNOR2_X1 i_71 (.A(add1_i[17]), .B(add2_i[17]), .ZN(n_54));
   XNOR2_X1 i_72 (.A(n_53), .B(n_54), .ZN(p_0[17]));
   INV_X1 i_73 (.A(add1_i[17]), .ZN(n_55));
   AOI22_X1 i_74 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(add2_i[17]), .ZN(n_56));
   XOR2_X1 i_75 (.A(add1_i[18]), .B(add2_i[18]), .Z(n_57));
   XNOR2_X1 i_76 (.A(n_56), .B(n_57), .ZN(p_0[18]));
   INV_X1 i_77 (.A(add2_i[18]), .ZN(n_58));
   OAI22_X1 i_78 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(add1_i[18]), .ZN(n_59));
   XNOR2_X1 i_79 (.A(add1_i[19]), .B(add2_i[19]), .ZN(n_60));
   XNOR2_X1 i_80 (.A(n_59), .B(n_60), .ZN(p_0[19]));
   INV_X1 i_81 (.A(add1_i[19]), .ZN(n_61));
   AOI22_X1 i_82 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(add2_i[19]), .ZN(n_62));
   XOR2_X1 i_83 (.A(add1_i[20]), .B(add2_i[20]), .Z(n_63));
   XNOR2_X1 i_84 (.A(n_62), .B(n_63), .ZN(p_0[20]));
   INV_X1 i_85 (.A(add2_i[20]), .ZN(n_64));
   OAI22_X1 i_86 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(add1_i[20]), .ZN(n_65));
   XNOR2_X1 i_87 (.A(add1_i[21]), .B(add2_i[21]), .ZN(n_66));
   XNOR2_X1 i_88 (.A(n_65), .B(n_66), .ZN(p_0[21]));
   INV_X1 i_89 (.A(add1_i[21]), .ZN(n_67));
   AOI22_X1 i_90 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(add2_i[21]), .ZN(n_68));
   XOR2_X1 i_91 (.A(add1_i[22]), .B(add2_i[22]), .Z(n_69));
   XNOR2_X1 i_92 (.A(n_68), .B(n_69), .ZN(p_0[22]));
   INV_X1 i_93 (.A(add2_i[22]), .ZN(n_70));
   OAI22_X1 i_94 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(add1_i[22]), .ZN(n_71));
   XNOR2_X1 i_95 (.A(add1_i[23]), .B(add2_i[23]), .ZN(n_72));
   XNOR2_X1 i_96 (.A(n_71), .B(n_72), .ZN(p_0[23]));
   INV_X1 i_97 (.A(add1_i[23]), .ZN(n_73));
   AOI22_X1 i_98 (.A1(n_71), .A2(n_72), .B1(n_73), .B2(add2_i[23]), .ZN(n_74));
   XOR2_X1 i_99 (.A(add1_i[24]), .B(add2_i[24]), .Z(n_75));
   XNOR2_X1 i_100 (.A(n_74), .B(n_75), .ZN(p_0[24]));
   INV_X1 i_101 (.A(add2_i[24]), .ZN(n_76));
   OAI22_X1 i_102 (.A1(n_74), .A2(n_75), .B1(n_76), .B2(add1_i[24]), .ZN(n_77));
   XNOR2_X1 i_103 (.A(add1_i[25]), .B(add2_i[25]), .ZN(n_78));
   XNOR2_X1 i_104 (.A(n_77), .B(n_78), .ZN(p_0[25]));
   INV_X1 i_105 (.A(add1_i[25]), .ZN(n_79));
   AOI22_X1 i_106 (.A1(n_77), .A2(n_78), .B1(n_79), .B2(add2_i[25]), .ZN(n_80));
   XOR2_X1 i_107 (.A(add1_i[26]), .B(add2_i[26]), .Z(n_81));
   XNOR2_X1 i_108 (.A(n_80), .B(n_81), .ZN(p_0[26]));
   INV_X1 i_109 (.A(add2_i[26]), .ZN(n_82));
   OAI22_X1 i_110 (.A1(n_80), .A2(n_81), .B1(n_82), .B2(add1_i[26]), .ZN(n_83));
   XOR2_X1 i_111 (.A(add2_i[27]), .B(add1_i[27]), .Z(n_84));
   XOR2_X1 i_112 (.A(n_83), .B(n_84), .Z(p_0[27]));
   INV_X1 i_113 (.A(n_83), .ZN(n_85));
   INV_X1 i_114 (.A(add2_i[27]), .ZN(n_86));
   OAI22_X1 i_115 (.A1(n_85), .A2(n_84), .B1(n_86), .B2(add1_i[27]), .ZN(p_0[28]));
endmodule

module datapath__0_55(add2_i, add1_i, p_0);
   input [27:0]add2_i;
   input [27:0]add1_i;
   output [28:0]p_0;

   HA_X1 i_0 (.A(add2_i[0]), .B(add1_i[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(add2_i[1]), .B(add1_i[1]), .CI(n_0), .CO(n_1), .S(p_0[1]));
   FA_X1 i_2 (.A(add2_i[2]), .B(add1_i[2]), .CI(n_1), .CO(n_2), .S(p_0[2]));
   FA_X1 i_3 (.A(add2_i[3]), .B(add1_i[3]), .CI(n_2), .CO(n_3), .S(p_0[3]));
   FA_X1 i_4 (.A(add2_i[4]), .B(add1_i[4]), .CI(n_3), .CO(n_4), .S(p_0[4]));
   FA_X1 i_5 (.A(add2_i[5]), .B(add1_i[5]), .CI(n_4), .CO(n_5), .S(p_0[5]));
   FA_X1 i_6 (.A(add2_i[6]), .B(add1_i[6]), .CI(n_5), .CO(n_6), .S(p_0[6]));
   FA_X1 i_7 (.A(add2_i[7]), .B(add1_i[7]), .CI(n_6), .CO(n_7), .S(p_0[7]));
   FA_X1 i_8 (.A(add2_i[8]), .B(add1_i[8]), .CI(n_7), .CO(n_8), .S(p_0[8]));
   FA_X1 i_9 (.A(add2_i[9]), .B(add1_i[9]), .CI(n_8), .CO(n_9), .S(p_0[9]));
   FA_X1 i_10 (.A(add2_i[10]), .B(add1_i[10]), .CI(n_9), .CO(n_10), .S(p_0[10]));
   FA_X1 i_11 (.A(add2_i[11]), .B(add1_i[11]), .CI(n_10), .CO(n_11), .S(p_0[11]));
   FA_X1 i_12 (.A(add2_i[12]), .B(add1_i[12]), .CI(n_11), .CO(n_12), .S(p_0[12]));
   FA_X1 i_13 (.A(add2_i[13]), .B(add1_i[13]), .CI(n_12), .CO(n_13), .S(p_0[13]));
   FA_X1 i_14 (.A(add2_i[14]), .B(add1_i[14]), .CI(n_13), .CO(n_14), .S(p_0[14]));
   FA_X1 i_15 (.A(add2_i[15]), .B(add1_i[15]), .CI(n_14), .CO(n_15), .S(p_0[15]));
   FA_X1 i_16 (.A(add2_i[16]), .B(add1_i[16]), .CI(n_15), .CO(n_16), .S(p_0[16]));
   FA_X1 i_17 (.A(add2_i[17]), .B(add1_i[17]), .CI(n_16), .CO(n_17), .S(p_0[17]));
   FA_X1 i_18 (.A(add2_i[18]), .B(add1_i[18]), .CI(n_17), .CO(n_18), .S(p_0[18]));
   FA_X1 i_19 (.A(add2_i[19]), .B(add1_i[19]), .CI(n_18), .CO(n_19), .S(p_0[19]));
   FA_X1 i_20 (.A(add2_i[20]), .B(add1_i[20]), .CI(n_19), .CO(n_20), .S(p_0[20]));
   FA_X1 i_21 (.A(add2_i[21]), .B(add1_i[21]), .CI(n_20), .CO(n_21), .S(p_0[21]));
   FA_X1 i_22 (.A(add2_i[22]), .B(add1_i[22]), .CI(n_21), .CO(n_22), .S(p_0[22]));
   FA_X1 i_23 (.A(add2_i[23]), .B(add1_i[23]), .CI(n_22), .CO(n_23), .S(p_0[23]));
   FA_X1 i_24 (.A(add2_i[24]), .B(add1_i[24]), .CI(n_23), .CO(n_24), .S(p_0[24]));
   FA_X1 i_25 (.A(add2_i[25]), .B(add1_i[25]), .CI(n_24), .CO(n_25), .S(p_0[25]));
   FA_X1 i_26 (.A(add2_i[26]), .B(add1_i[26]), .CI(n_25), .CO(n_26), .S(p_0[26]));
   FA_X1 i_27 (.A(add2_i[27]), .B(add1_i[27]), .CI(n_26), .CO(p_0[28]), .S(
      p_0[27]));
endmodule

module Adder(add1_i, add2_i, A_S, sum_o, carry_o);
   input [27:0]add1_i;
   input [27:0]add2_i;
   input A_S;
   output [27:0]sum_o;
   output carry_o;

   datapath__0_54 i_0 (.add1_i(add1_i), .p_0({n_28, n_27, n_26, n_25, n_24, n_23, 
      n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, 
      n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .add2_i(add2_i));
   datapath__0_55 i_1 (.add2_i(add2_i), .add1_i(add1_i), .p_0({n_57, n_56, n_55, 
      n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
      n_30, n_29}));
   MUX2_X1 i_2_0 (.A(n_29), .B(n_0), .S(A_S), .Z(sum_o[0]));
   MUX2_X1 i_2_1 (.A(n_30), .B(n_1), .S(A_S), .Z(sum_o[1]));
   MUX2_X1 i_2_2 (.A(n_31), .B(n_2), .S(A_S), .Z(sum_o[2]));
   MUX2_X1 i_2_3 (.A(n_32), .B(n_3), .S(A_S), .Z(sum_o[3]));
   MUX2_X1 i_2_4 (.A(n_33), .B(n_4), .S(A_S), .Z(sum_o[4]));
   MUX2_X1 i_2_5 (.A(n_34), .B(n_5), .S(A_S), .Z(sum_o[5]));
   MUX2_X1 i_2_6 (.A(n_35), .B(n_6), .S(A_S), .Z(sum_o[6]));
   MUX2_X1 i_2_7 (.A(n_36), .B(n_7), .S(A_S), .Z(sum_o[7]));
   MUX2_X1 i_2_8 (.A(n_37), .B(n_8), .S(A_S), .Z(sum_o[8]));
   MUX2_X1 i_2_9 (.A(n_38), .B(n_9), .S(A_S), .Z(sum_o[9]));
   MUX2_X1 i_2_10 (.A(n_39), .B(n_10), .S(A_S), .Z(sum_o[10]));
   MUX2_X1 i_2_11 (.A(n_40), .B(n_11), .S(A_S), .Z(sum_o[11]));
   MUX2_X1 i_2_12 (.A(n_41), .B(n_12), .S(A_S), .Z(sum_o[12]));
   MUX2_X1 i_2_13 (.A(n_42), .B(n_13), .S(A_S), .Z(sum_o[13]));
   MUX2_X1 i_2_14 (.A(n_43), .B(n_14), .S(A_S), .Z(sum_o[14]));
   MUX2_X1 i_2_15 (.A(n_44), .B(n_15), .S(A_S), .Z(sum_o[15]));
   MUX2_X1 i_2_16 (.A(n_45), .B(n_16), .S(A_S), .Z(sum_o[16]));
   MUX2_X1 i_2_17 (.A(n_46), .B(n_17), .S(A_S), .Z(sum_o[17]));
   MUX2_X1 i_2_18 (.A(n_47), .B(n_18), .S(A_S), .Z(sum_o[18]));
   MUX2_X1 i_2_19 (.A(n_48), .B(n_19), .S(A_S), .Z(sum_o[19]));
   MUX2_X1 i_2_20 (.A(n_49), .B(n_20), .S(A_S), .Z(sum_o[20]));
   MUX2_X1 i_2_21 (.A(n_50), .B(n_21), .S(A_S), .Z(sum_o[21]));
   MUX2_X1 i_2_22 (.A(n_51), .B(n_22), .S(A_S), .Z(sum_o[22]));
   MUX2_X1 i_2_23 (.A(n_52), .B(n_23), .S(A_S), .Z(sum_o[23]));
   MUX2_X1 i_2_24 (.A(n_53), .B(n_24), .S(A_S), .Z(sum_o[24]));
   MUX2_X1 i_2_25 (.A(n_54), .B(n_25), .S(A_S), .Z(sum_o[25]));
   MUX2_X1 i_2_26 (.A(n_55), .B(n_26), .S(A_S), .Z(sum_o[26]));
   MUX2_X1 i_2_27 (.A(n_56), .B(n_27), .S(A_S), .Z(sum_o[27]));
   MUX2_X1 i_2_28 (.A(n_57), .B(n_28), .S(A_S), .Z(carry_o));
endmodule

module datapath__0_58(p_0, p_1);
   input [27:0]p_0;
   output [27:0]p_1;

   HA_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_1 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_2 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_3 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
   HA_X1 i_4 (.A(p_0[5]), .B(n_3), .CO(n_4), .S(p_1[5]));
   HA_X1 i_5 (.A(p_0[6]), .B(n_4), .CO(n_5), .S(p_1[6]));
   HA_X1 i_6 (.A(p_0[7]), .B(n_5), .CO(n_6), .S(p_1[7]));
   HA_X1 i_7 (.A(p_0[8]), .B(n_6), .CO(n_7), .S(p_1[8]));
   HA_X1 i_8 (.A(p_0[9]), .B(n_7), .CO(n_8), .S(p_1[9]));
   HA_X1 i_9 (.A(p_0[10]), .B(n_8), .CO(n_9), .S(p_1[10]));
   HA_X1 i_10 (.A(p_0[11]), .B(n_9), .CO(n_10), .S(p_1[11]));
   HA_X1 i_11 (.A(p_0[12]), .B(n_10), .CO(n_11), .S(p_1[12]));
   HA_X1 i_12 (.A(p_0[13]), .B(n_11), .CO(n_12), .S(p_1[13]));
   HA_X1 i_13 (.A(p_0[14]), .B(n_12), .CO(n_13), .S(p_1[14]));
   HA_X1 i_14 (.A(p_0[15]), .B(n_13), .CO(n_14), .S(p_1[15]));
   HA_X1 i_15 (.A(p_0[16]), .B(n_14), .CO(n_15), .S(p_1[16]));
   HA_X1 i_16 (.A(p_0[17]), .B(n_15), .CO(n_16), .S(p_1[17]));
   HA_X1 i_17 (.A(p_0[18]), .B(n_16), .CO(n_17), .S(p_1[18]));
   HA_X1 i_18 (.A(p_0[19]), .B(n_17), .CO(n_18), .S(p_1[19]));
   HA_X1 i_19 (.A(p_0[20]), .B(n_18), .CO(n_19), .S(p_1[20]));
   HA_X1 i_20 (.A(p_0[21]), .B(n_19), .CO(n_20), .S(p_1[21]));
   HA_X1 i_21 (.A(p_0[22]), .B(n_20), .CO(n_21), .S(p_1[22]));
   HA_X1 i_22 (.A(p_0[23]), .B(n_21), .CO(n_22), .S(p_1[23]));
   HA_X1 i_23 (.A(p_0[24]), .B(n_22), .CO(n_23), .S(p_1[24]));
   HA_X1 i_24 (.A(p_0[25]), .B(n_23), .CO(n_24), .S(p_1[25]));
   HA_X1 i_25 (.A(p_0[26]), .B(n_24), .CO(n_25), .S(p_1[26]));
   XOR2_X1 i_26 (.A(p_0[27]), .B(n_25), .Z(p_1[27]));
endmodule

module block_adder(SA, SB, Comp, A, B, A_S, MS, CO, SO);
   input SA;
   input SB;
   input Comp;
   input [27:0]A;
   input [27:0]B;
   input A_S;
   output [27:0]MS;
   output CO;
   output SO;

   wire AS_aux;
   wire [27:0]Bb_aux;
   wire [27:0]Aa_aux;
   wire CO_aux;
   wire [27:0]MS_aux;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   signout so (.SA(SA), .SB(SB), .Comp(Comp), .A({A[27], A[26], A[25], A[24], 
      A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], uc_0, uc_1, 
      uc_2, uc_3}), .B(B), .A_S(A_S), .Aa(Aa_aux), .Bb(Bb_aux), .AS(AS_aux), 
      .SO(SO));
   Adder add (.add1_i(Aa_aux), .add2_i(Bb_aux), .A_S(AS_aux), .sum_o({MS_aux[27], 
      MS_aux[26], MS_aux[25], MS_aux[24], MS_aux[23], MS_aux[22], MS_aux[21], 
      MS_aux[20], MS_aux[19], MS_aux[18], MS_aux[17], MS_aux[16], MS_aux[15], 
      MS_aux[14], MS_aux[13], MS_aux[12], MS_aux[11], MS_aux[10], MS_aux[9], 
      MS_aux[8], MS_aux[7], MS_aux[6], MS_aux[5], MS_aux[4], MS_aux[3], 
      MS_aux[2], MS_aux[1], MS[0]}), .carry_o(CO_aux));
   datapath__0_58 i_1 (.p_0({n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, 
      n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, 
      n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27}), .p_1({n_26, n_25, n_24, 
      n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, 
      n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_4}));
   AND2_X1 i_0_0 (.A1(n_0_0), .A2(CO_aux), .ZN(CO));
   XNOR2_X1 i_0_1 (.A(SA), .B(n_0_1), .ZN(n_0_0));
   XOR2_X1 i_0_2 (.A(A_S), .B(SB), .Z(n_0_1));
   MUX2_X1 i_0_3 (.A(n_0), .B(MS_aux[1]), .S(n_0_2), .Z(MS[1]));
   MUX2_X1 i_0_4 (.A(n_1), .B(MS_aux[2]), .S(n_0_2), .Z(MS[2]));
   MUX2_X1 i_0_5 (.A(n_2), .B(MS_aux[3]), .S(n_0_2), .Z(MS[3]));
   MUX2_X1 i_0_6 (.A(n_3), .B(MS_aux[4]), .S(n_0_2), .Z(MS[4]));
   MUX2_X1 i_0_7 (.A(n_4), .B(MS_aux[5]), .S(n_0_2), .Z(MS[5]));
   MUX2_X1 i_0_8 (.A(n_5), .B(MS_aux[6]), .S(n_0_2), .Z(MS[6]));
   MUX2_X1 i_0_9 (.A(n_6), .B(MS_aux[7]), .S(n_0_2), .Z(MS[7]));
   MUX2_X1 i_0_10 (.A(n_7), .B(MS_aux[8]), .S(n_0_2), .Z(MS[8]));
   MUX2_X1 i_0_11 (.A(n_8), .B(MS_aux[9]), .S(n_0_2), .Z(MS[9]));
   MUX2_X1 i_0_12 (.A(n_9), .B(MS_aux[10]), .S(n_0_2), .Z(MS[10]));
   MUX2_X1 i_0_13 (.A(n_10), .B(MS_aux[11]), .S(n_0_2), .Z(MS[11]));
   MUX2_X1 i_0_14 (.A(n_11), .B(MS_aux[12]), .S(n_0_2), .Z(MS[12]));
   MUX2_X1 i_0_15 (.A(n_12), .B(MS_aux[13]), .S(n_0_2), .Z(MS[13]));
   MUX2_X1 i_0_16 (.A(n_13), .B(MS_aux[14]), .S(n_0_2), .Z(MS[14]));
   MUX2_X1 i_0_17 (.A(n_14), .B(MS_aux[15]), .S(n_0_2), .Z(MS[15]));
   MUX2_X1 i_0_18 (.A(n_15), .B(MS_aux[16]), .S(n_0_2), .Z(MS[16]));
   MUX2_X1 i_0_19 (.A(n_16), .B(MS_aux[17]), .S(n_0_2), .Z(MS[17]));
   MUX2_X1 i_0_20 (.A(n_17), .B(MS_aux[18]), .S(n_0_2), .Z(MS[18]));
   MUX2_X1 i_0_21 (.A(n_18), .B(MS_aux[19]), .S(n_0_2), .Z(MS[19]));
   MUX2_X1 i_0_22 (.A(n_19), .B(MS_aux[20]), .S(n_0_2), .Z(MS[20]));
   MUX2_X1 i_0_23 (.A(n_20), .B(MS_aux[21]), .S(n_0_2), .Z(MS[21]));
   MUX2_X1 i_0_24 (.A(n_21), .B(MS_aux[22]), .S(n_0_2), .Z(MS[22]));
   MUX2_X1 i_0_25 (.A(n_22), .B(MS_aux[23]), .S(n_0_2), .Z(MS[23]));
   MUX2_X1 i_0_26 (.A(n_23), .B(MS_aux[24]), .S(n_0_2), .Z(MS[24]));
   MUX2_X1 i_0_27 (.A(n_24), .B(MS_aux[25]), .S(n_0_2), .Z(MS[25]));
   MUX2_X1 i_0_28 (.A(n_25), .B(MS_aux[26]), .S(n_0_2), .Z(MS[26]));
   MUX2_X1 i_0_29 (.A(n_26), .B(MS_aux[27]), .S(n_0_2), .Z(MS[27]));
   NAND2_X1 i_0_30 (.A1(SO), .A2(AS_aux), .ZN(n_0_2));
   INV_X1 i_0_31 (.A(MS[0]), .ZN(n_27));
   INV_X1 i_0_32 (.A(MS_aux[1]), .ZN(n_28));
   INV_X1 i_0_33 (.A(MS_aux[2]), .ZN(n_29));
   INV_X1 i_0_34 (.A(MS_aux[3]), .ZN(n_30));
   INV_X1 i_0_35 (.A(MS_aux[4]), .ZN(n_31));
   INV_X1 i_0_36 (.A(MS_aux[5]), .ZN(n_32));
   INV_X1 i_0_37 (.A(MS_aux[6]), .ZN(n_33));
   INV_X1 i_0_38 (.A(MS_aux[7]), .ZN(n_34));
   INV_X1 i_0_39 (.A(MS_aux[8]), .ZN(n_35));
   INV_X1 i_0_40 (.A(MS_aux[9]), .ZN(n_36));
   INV_X1 i_0_41 (.A(MS_aux[10]), .ZN(n_37));
   INV_X1 i_0_42 (.A(MS_aux[11]), .ZN(n_38));
   INV_X1 i_0_43 (.A(MS_aux[12]), .ZN(n_39));
   INV_X1 i_0_44 (.A(MS_aux[13]), .ZN(n_40));
   INV_X1 i_0_45 (.A(MS_aux[14]), .ZN(n_41));
   INV_X1 i_0_46 (.A(MS_aux[15]), .ZN(n_42));
   INV_X1 i_0_47 (.A(MS_aux[16]), .ZN(n_43));
   INV_X1 i_0_48 (.A(MS_aux[17]), .ZN(n_44));
   INV_X1 i_0_49 (.A(MS_aux[18]), .ZN(n_45));
   INV_X1 i_0_50 (.A(MS_aux[19]), .ZN(n_46));
   INV_X1 i_0_51 (.A(MS_aux[20]), .ZN(n_47));
   INV_X1 i_0_52 (.A(MS_aux[21]), .ZN(n_48));
   INV_X1 i_0_53 (.A(MS_aux[22]), .ZN(n_49));
   INV_X1 i_0_54 (.A(MS_aux[23]), .ZN(n_50));
   INV_X1 i_0_55 (.A(MS_aux[24]), .ZN(n_51));
   INV_X1 i_0_56 (.A(MS_aux[25]), .ZN(n_52));
   INV_X1 i_0_57 (.A(MS_aux[26]), .ZN(n_53));
   INV_X1 i_0_58 (.A(MS_aux[27]), .ZN(n_54));
endmodule

module zero_counter(M, Zcount);
   input [27:0]M;
   output [4:0]Zcount;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;

   OR4_X1 i_0_0 (.A1(n_0_13), .A2(n_0_4), .A3(n_0_1), .A4(n_0_0), .ZN(Zcount[0]));
   NOR3_X1 i_0_1 (.A1(n_0_29), .A2(n_0_2), .A3(M[7]), .ZN(n_0_0));
   NOR3_X1 i_0_2 (.A1(n_0_32), .A2(n_0_3), .A3(M[11]), .ZN(n_0_1));
   AOI21_X1 i_0_3 (.A(M[6]), .B1(n_0_42), .B2(M[4]), .ZN(n_0_2));
   AOI21_X1 i_0_4 (.A(M[10]), .B1(n_0_43), .B2(M[8]), .ZN(n_0_3));
   NOR2_X1 i_0_5 (.A1(Zcount[4]), .A2(n_0_5), .ZN(n_0_4));
   OAI21_X1 i_0_6 (.A(n_0_9), .B1(n_0_6), .B2(n_0_36), .ZN(n_0_5));
   NOR2_X1 i_0_7 (.A1(M[17]), .A2(n_0_7), .ZN(n_0_6));
   NOR2_X1 i_0_8 (.A1(M[16]), .A2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(M[15]), .B1(n_0_44), .B2(M[13]), .ZN(n_0_8));
   OAI22_X1 i_0_10 (.A1(n_0_10), .A2(M[27]), .B1(n_0_37), .B2(M[19]), .ZN(n_0_9));
   OAI211_X1 i_0_11 (.A(n_0_37), .B(n_0_11), .C1(M[26]), .C2(n_0_46), .ZN(n_0_10));
   OAI21_X1 i_0_12 (.A(n_0_40), .B1(n_0_12), .B2(M[23]), .ZN(n_0_11));
   NOR2_X1 i_0_13 (.A1(n_0_45), .A2(M[22]), .ZN(n_0_12));
   NOR3_X1 i_0_14 (.A1(n_0_27), .A2(n_0_14), .A3(M[3]), .ZN(n_0_13));
   AOI21_X1 i_0_15 (.A(M[2]), .B1(n_0_41), .B2(M[0]), .ZN(n_0_14));
   OAI21_X1 i_0_16 (.A(n_0_15), .B1(n_0_25), .B2(n_0_26), .ZN(Zcount[1]));
   OAI211_X1 i_0_17 (.A(n_0_27), .B(n_0_17), .C1(n_0_16), .C2(n_0_32), .ZN(
      n_0_15));
   AOI211_X1 i_0_18 (.A(M[11]), .B(M[10]), .C1(n_0_28), .C2(n_0_31), .ZN(n_0_16));
   OAI21_X1 i_0_19 (.A(n_0_18), .B1(n_0_36), .B2(n_0_21), .ZN(n_0_17));
   NAND2_X1 i_0_20 (.A1(n_0_19), .A2(n_0_37), .ZN(n_0_18));
   NOR3_X1 i_0_21 (.A1(M[27]), .A2(M[26]), .A3(n_0_20), .ZN(n_0_19));
   NOR3_X1 i_0_22 (.A1(M[25]), .A2(M[24]), .A3(n_0_39), .ZN(n_0_20));
   NOR3_X1 i_0_23 (.A1(M[17]), .A2(M[16]), .A3(n_0_34), .ZN(n_0_21));
   INV_X1 i_0_24 (.A(n_0_22), .ZN(Zcount[2]));
   AOI21_X1 i_0_25 (.A(n_0_25), .B1(n_0_23), .B2(n_0_27), .ZN(n_0_22));
   OAI21_X1 i_0_26 (.A(n_0_29), .B1(n_0_24), .B2(Zcount[4]), .ZN(n_0_23));
   AOI21_X1 i_0_27 (.A(n_0_35), .B1(n_0_37), .B2(n_0_40), .ZN(n_0_24));
   NOR3_X1 i_0_28 (.A1(n_0_26), .A2(M[0]), .A3(M[1]), .ZN(n_0_25));
   OR3_X1 i_0_29 (.A1(n_0_27), .A2(M[2]), .A3(M[3]), .ZN(n_0_26));
   OAI21_X1 i_0_30 (.A(n_0_27), .B1(Zcount[4]), .B2(n_0_37), .ZN(Zcount[3]));
   OR4_X1 i_0_31 (.A1(n_0_29), .A2(n_0_28), .A3(M[5]), .A4(M[4]), .ZN(n_0_27));
   OR2_X1 i_0_32 (.A1(M[7]), .A2(M[6]), .ZN(n_0_28));
   NAND3_X1 i_0_33 (.A1(Zcount[4]), .A2(n_0_31), .A3(n_0_30), .ZN(n_0_29));
   NOR2_X1 i_0_34 (.A1(M[11]), .A2(M[10]), .ZN(n_0_30));
   NOR2_X1 i_0_35 (.A1(M[9]), .A2(M[8]), .ZN(n_0_31));
   INV_X1 i_0_36 (.A(Zcount[4]), .ZN(n_0_32));
   AND3_X1 i_0_37 (.A1(n_0_35), .A2(n_0_34), .A3(n_0_33), .ZN(Zcount[4]));
   NOR2_X1 i_0_38 (.A1(M[13]), .A2(M[12]), .ZN(n_0_33));
   NOR2_X1 i_0_39 (.A1(M[15]), .A2(M[14]), .ZN(n_0_34));
   NOR3_X1 i_0_40 (.A1(n_0_36), .A2(M[16]), .A3(M[17]), .ZN(n_0_35));
   OR3_X1 i_0_41 (.A1(n_0_37), .A2(M[18]), .A3(M[19]), .ZN(n_0_36));
   NAND3_X1 i_0_42 (.A1(n_0_40), .A2(n_0_39), .A3(n_0_38), .ZN(n_0_37));
   NOR2_X1 i_0_43 (.A1(M[21]), .A2(M[20]), .ZN(n_0_38));
   NOR2_X1 i_0_44 (.A1(M[23]), .A2(M[22]), .ZN(n_0_39));
   NOR4_X1 i_0_45 (.A1(M[27]), .A2(M[26]), .A3(M[25]), .A4(M[24]), .ZN(n_0_40));
   INV_X1 i_0_46 (.A(M[1]), .ZN(n_0_41));
   INV_X1 i_0_47 (.A(M[5]), .ZN(n_0_42));
   INV_X1 i_0_48 (.A(M[9]), .ZN(n_0_43));
   INV_X1 i_0_49 (.A(M[14]), .ZN(n_0_44));
   INV_X1 i_0_50 (.A(M[21]), .ZN(n_0_45));
   INV_X1 i_0_51 (.A(M[25]), .ZN(n_0_46));
endmodule

module exponent(ES, Co, Zcount_aux, shift, E);
   input [7:0]ES;
   input Co;
   input [4:0]Zcount_aux;
   output [4:0]shift;
   output [7:0]E;

   wire n_0_0;
   wire n_0_17;
   wire n_0_4;
   wire n_0_18;
   wire n_0_7;
   wire n_0_19;
   wire n_0_10;
   wire n_0_20;
   wire n_0_13;
   wire n_0_21;
   wire n_0_16;
   wire n_0_22;
   wire n_0_11;
   wire n_0_8;
   wire n_0_5;
   wire n_0_2;
   wire n_0_23;
   wire n_0_24;
   wire n_0_15;
   wire n_0_25;
   wire n_0_1;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_12;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_6;
   wire n_0_9;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_3;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_14;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;

   FA_X1 i_0_0 (.A(n_0_1), .B(n_0_2), .CI(n_0_15), .CO(n_0_17), .S(n_0_0));
   FA_X1 i_0_1 (.A(n_0_3), .B(n_0_5), .CI(n_0_17), .CO(n_0_18), .S(n_0_4));
   FA_X1 i_0_2 (.A(n_0_6), .B(n_0_8), .CI(n_0_18), .CO(n_0_19), .S(n_0_7));
   FA_X1 i_0_3 (.A(n_0_9), .B(n_0_11), .CI(n_0_19), .CO(n_0_20), .S(n_0_10));
   FA_X1 i_0_4 (.A(n_0_12), .B(n_0_14), .CI(n_0_20), .CO(n_0_21), .S(n_0_13));
   FA_X1 i_0_5 (.A(ES[6]), .B(n_0_14), .CI(n_0_21), .CO(n_0_22), .S(n_0_16));
   NOR2_X1 i_0_6 (.A1(n_0_44), .A2(n_0_12), .ZN(n_0_11));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_43), .ZN(n_0_8));
   NOR2_X1 i_0_8 (.A1(n_0_47), .A2(n_0_6), .ZN(n_0_5));
   NOR2_X1 i_0_9 (.A1(n_0_3), .A2(n_0_48), .ZN(n_0_2));
   AOI21_X1 i_0_10 (.A(n_0_23), .B1(n_0_24), .B2(n_0_29), .ZN(E[0]));
   NAND2_X1 i_0_11 (.A1(n_0_40), .A2(n_0_34), .ZN(n_0_23));
   XNOR2_X1 i_0_12 (.A(Zcount_aux[0]), .B(n_0_25), .ZN(n_0_24));
   NOR2_X1 i_0_13 (.A1(Zcount_aux[0]), .A2(n_0_25), .ZN(n_0_15));
   XOR2_X1 i_0_14 (.A(ES[0]), .B(Co), .Z(n_0_25));
   OR2_X1 i_0_15 (.A1(ES[0]), .A2(Co), .ZN(n_0_1));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(n_0_28), .ZN(E[1]));
   AND2_X1 i_0_17 (.A1(n_0_4), .A2(n_0_28), .ZN(E[2]));
   AND2_X1 i_0_18 (.A1(n_0_7), .A2(n_0_28), .ZN(E[3]));
   AND2_X1 i_0_19 (.A1(n_0_10), .A2(n_0_28), .ZN(E[4]));
   AND2_X1 i_0_20 (.A1(n_0_13), .A2(n_0_28), .ZN(E[5]));
   AND2_X1 i_0_21 (.A1(n_0_16), .A2(n_0_28), .ZN(E[6]));
   AND2_X1 i_0_22 (.A1(n_0_28), .A2(n_0_26), .ZN(E[7]));
   XNOR2_X1 i_0_23 (.A(n_0_22), .B(n_0_27), .ZN(n_0_26));
   XNOR2_X1 i_0_24 (.A(ES[7]), .B(n_0_14), .ZN(n_0_27));
   AND2_X1 i_0_25 (.A1(n_0_34), .A2(n_0_29), .ZN(n_0_28));
   OAI21_X1 i_0_26 (.A(n_0_50), .B1(n_0_44), .B2(n_0_30), .ZN(n_0_29));
   NOR3_X1 i_0_27 (.A1(n_0_9), .A2(n_0_12), .A3(n_0_31), .ZN(n_0_30));
   NOR3_X1 i_0_28 (.A1(n_0_47), .A2(n_0_43), .A3(n_0_32), .ZN(n_0_31));
   AOI211_X1 i_0_29 (.A(n_0_3), .B(n_0_6), .C1(n_0_33), .C2(ES[0]), .ZN(n_0_32));
   NOR2_X1 i_0_30 (.A1(Zcount_aux[0]), .A2(n_0_48), .ZN(n_0_33));
   NAND3_X1 i_0_31 (.A1(Zcount_aux[4]), .A2(Zcount_aux[3]), .A3(n_0_35), 
      .ZN(n_0_34));
   NOR3_X1 i_0_32 (.A1(n_0_55), .A2(Zcount_aux[1]), .A3(Zcount_aux[0]), .ZN(
      n_0_35));
   AOI21_X1 i_0_33 (.A(n_0_36), .B1(n_0_40), .B2(n_0_54), .ZN(shift[0]));
   NOR2_X1 i_0_34 (.A1(n_0_40), .A2(ES[0]), .ZN(n_0_36));
   OAI21_X1 i_0_35 (.A(n_0_37), .B1(n_0_40), .B2(n_0_51), .ZN(shift[1]));
   NAND2_X1 i_0_36 (.A1(n_0_40), .A2(Zcount_aux[1]), .ZN(n_0_37));
   AOI21_X1 i_0_37 (.A(n_0_38), .B1(n_0_40), .B2(n_0_55), .ZN(shift[2]));
   NOR2_X1 i_0_38 (.A1(n_0_40), .A2(ES[2]), .ZN(n_0_38));
   OAI21_X1 i_0_39 (.A(n_0_39), .B1(n_0_40), .B2(n_0_52), .ZN(shift[3]));
   NAND2_X1 i_0_40 (.A1(n_0_40), .A2(Zcount_aux[3]), .ZN(n_0_39));
   NAND2_X1 i_0_41 (.A1(n_0_50), .A2(n_0_41), .ZN(n_0_40));
   NOR2_X1 i_0_42 (.A1(n_0_42), .A2(n_0_12), .ZN(n_0_41));
   NOR2_X1 i_0_43 (.A1(n_0_53), .A2(Zcount_aux[4]), .ZN(n_0_12));
   NOR3_X1 i_0_44 (.A1(n_0_45), .A2(n_0_44), .A3(n_0_43), .ZN(n_0_42));
   AND2_X1 i_0_45 (.A1(n_0_52), .A2(Zcount_aux[3]), .ZN(n_0_43));
   NOR2_X1 i_0_46 (.A1(n_0_56), .A2(ES[4]), .ZN(n_0_44));
   NOR3_X1 i_0_47 (.A1(n_0_46), .A2(n_0_9), .A3(n_0_6), .ZN(n_0_45));
   AND2_X1 i_0_48 (.A1(n_0_55), .A2(ES[2]), .ZN(n_0_6));
   NOR2_X1 i_0_49 (.A1(n_0_52), .A2(Zcount_aux[3]), .ZN(n_0_9));
   NOR3_X1 i_0_50 (.A1(n_0_49), .A2(n_0_48), .A3(n_0_47), .ZN(n_0_46));
   NOR2_X1 i_0_51 (.A1(n_0_55), .A2(ES[2]), .ZN(n_0_47));
   AND2_X1 i_0_52 (.A1(n_0_51), .A2(Zcount_aux[1]), .ZN(n_0_48));
   NOR3_X1 i_0_53 (.A1(n_0_3), .A2(n_0_54), .A3(ES[0]), .ZN(n_0_49));
   NOR2_X1 i_0_54 (.A1(n_0_51), .A2(Zcount_aux[1]), .ZN(n_0_3));
   AOI21_X1 i_0_55 (.A(n_0_56), .B1(n_0_50), .B2(n_0_53), .ZN(shift[4]));
   NOR3_X1 i_0_56 (.A1(ES[7]), .A2(ES[6]), .A3(ES[5]), .ZN(n_0_50));
   INV_X1 i_0_57 (.A(ES[1]), .ZN(n_0_51));
   INV_X1 i_0_58 (.A(ES[3]), .ZN(n_0_52));
   INV_X1 i_0_59 (.A(ES[4]), .ZN(n_0_53));
   INV_X1 i_0_60 (.A(ES[5]), .ZN(n_0_14));
   INV_X1 i_0_61 (.A(Zcount_aux[0]), .ZN(n_0_54));
   INV_X1 i_0_62 (.A(Zcount_aux[2]), .ZN(n_0_55));
   INV_X1 i_0_63 (.A(Zcount_aux[4]), .ZN(n_0_56));
endmodule

module mux2X1__0_77(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_79(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_81(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_83(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_85(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_87(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_89(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_91(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_93(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_95(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_97(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_99(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_101(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_103(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_105(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_107(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_109(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_111(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_113(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_115(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_117(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_119(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_121(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_123(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_125(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_127(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_129(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_131(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_133(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_135(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_137(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_139(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_141(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_143(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_145(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_147(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_149(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_151(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_153(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_155(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_157(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_159(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_161(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_163(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_165(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_167(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_169(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_171(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_173(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_175(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_177(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_179(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_181(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_183(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_185(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_187(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_189(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_191(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_193(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_195(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_197(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_199(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_201(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_203(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_205(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_207(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_209(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_211(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_213(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_215(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_217(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_219(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_221(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_223(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_225(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_227(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_229(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_231(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_233(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_235(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_237(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_239(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_241(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_243(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_245(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_247(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_249(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_251(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_253(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_255(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_257(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_259(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_261(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_263(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_265(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_267(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_269(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_271(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_273(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_275(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_277(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_279(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_281(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_283(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_285(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_287(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_289(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_291(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_293(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_295(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_297(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_299(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_301(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   wire n_0_0;

   INV_X1 i_0_0 (.A(in1), .ZN(n_0_0));
   NOR2_X1 i_0_1 (.A1(n_0_0), .A2(sel), .ZN(out));
endmodule

module mux2X1__0_303(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_305(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_307(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_309(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_311(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_313(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_315(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_317(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_319(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_321(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_323(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_325(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_327(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_329(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_331(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_333(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_335(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_337(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_339(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_341(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_343(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_345(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_347(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_349(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_351(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1__0_353(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module mux2X1(in0, in1, sel, out);
   input in0;
   input in1;
   input sel;
   output out;

   MUX2_X1 i_0_0 (.A(in1), .B(in0), .S(sel), .Z(out));
endmodule

module n_shift(shft, in, out);
   input [4:0]shft;
   input [27:0]in;
   output [27:0]out;

   wire [27:0]z4;
   wire [27:0]z3;
   wire [27:0]z2;
   wire [27:0]z1;

   mux2X1__0_77 genblk1_0_m9 (.in0(), .in1(z4[0]), .sel(shft[4]), .out(out[0]));
   mux2X1__0_79 genblk1_1_m9 (.in0(), .in1(z4[1]), .sel(shft[4]), .out(out[1]));
   mux2X1__0_81 genblk1_2_m9 (.in0(), .in1(z4[2]), .sel(shft[4]), .out(out[2]));
   mux2X1__0_83 genblk1_3_m9 (.in0(), .in1(z4[3]), .sel(shft[4]), .out(out[3]));
   mux2X1__0_85 genblk1_4_m9 (.in0(), .in1(z4[4]), .sel(shft[4]), .out(out[4]));
   mux2X1__0_87 genblk1_5_m9 (.in0(), .in1(z4[5]), .sel(shft[4]), .out(out[5]));
   mux2X1__0_89 genblk1_6_m9 (.in0(), .in1(z4[6]), .sel(shft[4]), .out(out[6]));
   mux2X1__0_91 genblk1_7_m9 (.in0(), .in1(z4[7]), .sel(shft[4]), .out(out[7]));
   mux2X1__0_93 genblk1_8_m9 (.in0(), .in1(z4[8]), .sel(shft[4]), .out(out[8]));
   mux2X1__0_95 genblk1_9_m9 (.in0(), .in1(z4[9]), .sel(shft[4]), .out(out[9]));
   mux2X1__0_97 genblk1_10_m9 (.in0(), .in1(z4[10]), .sel(shft[4]), .out(out[10]));
   mux2X1__0_99 genblk1_11_m9 (.in0(), .in1(z4[11]), .sel(shft[4]), .out(out[11]));
   mux2X1__0_101 genblk1_12_m9 (.in0(), .in1(z4[12]), .sel(shft[4]), .out(
      out[12]));
   mux2X1__0_103 genblk1_13_m9 (.in0(), .in1(z4[13]), .sel(shft[4]), .out(
      out[13]));
   mux2X1__0_105 genblk1_14_m9 (.in0(), .in1(z4[14]), .sel(shft[4]), .out(
      out[14]));
   mux2X1__0_107 genblk1_15_m9 (.in0(), .in1(z4[15]), .sel(shft[4]), .out(
      out[15]));
   mux2X1__0_109 genblk1_16_m10 (.in0(z4[0]), .in1(z4[16]), .sel(shft[4]), 
      .out(out[16]));
   mux2X1__0_111 genblk1_17_m10 (.in0(z4[1]), .in1(z4[17]), .sel(shft[4]), 
      .out(out[17]));
   mux2X1__0_113 genblk1_18_m10 (.in0(z4[2]), .in1(z4[18]), .sel(shft[4]), 
      .out(out[18]));
   mux2X1__0_115 genblk1_19_m10 (.in0(z4[3]), .in1(z4[19]), .sel(shft[4]), 
      .out(out[19]));
   mux2X1__0_117 genblk1_20_m10 (.in0(z4[4]), .in1(z4[20]), .sel(shft[4]), 
      .out(out[20]));
   mux2X1__0_119 genblk1_21_m10 (.in0(z4[5]), .in1(z4[21]), .sel(shft[4]), 
      .out(out[21]));
   mux2X1__0_121 genblk1_22_m10 (.in0(z4[6]), .in1(z4[22]), .sel(shft[4]), 
      .out(out[22]));
   mux2X1__0_123 genblk1_23_m10 (.in0(z4[7]), .in1(z4[23]), .sel(shft[4]), 
      .out(out[23]));
   mux2X1__0_125 genblk1_24_m10 (.in0(z4[8]), .in1(z4[24]), .sel(shft[4]), 
      .out(out[24]));
   mux2X1__0_127 genblk1_25_m10 (.in0(z4[9]), .in1(z4[25]), .sel(shft[4]), 
      .out(out[25]));
   mux2X1__0_129 genblk1_26_m10 (.in0(z4[10]), .in1(z4[26]), .sel(shft[4]), 
      .out(out[26]));
   mux2X1__0_131 genblk1_27_m10 (.in0(z4[11]), .in1(z4[27]), .sel(shft[4]), 
      .out(out[27]));
   mux2X1__0_133 genblk1_0_m7 (.in0(), .in1(z3[0]), .sel(shft[3]), .out(z4[0]));
   mux2X1__0_135 genblk1_1_m7 (.in0(), .in1(z3[1]), .sel(shft[3]), .out(z4[1]));
   mux2X1__0_137 genblk1_2_m7 (.in0(), .in1(z3[2]), .sel(shft[3]), .out(z4[2]));
   mux2X1__0_139 genblk1_3_m7 (.in0(), .in1(z3[3]), .sel(shft[3]), .out(z4[3]));
   mux2X1__0_141 genblk1_4_m7 (.in0(), .in1(z3[4]), .sel(shft[3]), .out(z4[4]));
   mux2X1__0_143 genblk1_5_m7 (.in0(), .in1(z3[5]), .sel(shft[3]), .out(z4[5]));
   mux2X1__0_145 genblk1_6_m7 (.in0(), .in1(z3[6]), .sel(shft[3]), .out(z4[6]));
   mux2X1__0_147 genblk1_7_m7 (.in0(), .in1(z3[7]), .sel(shft[3]), .out(z4[7]));
   mux2X1__0_149 genblk1_8_m8 (.in0(z3[0]), .in1(z3[8]), .sel(shft[3]), .out(
      z4[8]));
   mux2X1__0_151 genblk1_9_m8 (.in0(z3[1]), .in1(z3[9]), .sel(shft[3]), .out(
      z4[9]));
   mux2X1__0_153 genblk1_10_m8 (.in0(z3[2]), .in1(z3[10]), .sel(shft[3]), 
      .out(z4[10]));
   mux2X1__0_155 genblk1_11_m8 (.in0(z3[3]), .in1(z3[11]), .sel(shft[3]), 
      .out(z4[11]));
   mux2X1__0_157 genblk1_12_m8 (.in0(z3[4]), .in1(z3[12]), .sel(shft[3]), 
      .out(z4[12]));
   mux2X1__0_159 genblk1_13_m8 (.in0(z3[5]), .in1(z3[13]), .sel(shft[3]), 
      .out(z4[13]));
   mux2X1__0_161 genblk1_14_m8 (.in0(z3[6]), .in1(z3[14]), .sel(shft[3]), 
      .out(z4[14]));
   mux2X1__0_163 genblk1_15_m8 (.in0(z3[7]), .in1(z3[15]), .sel(shft[3]), 
      .out(z4[15]));
   mux2X1__0_165 genblk1_16_m8 (.in0(z3[8]), .in1(z3[16]), .sel(shft[3]), 
      .out(z4[16]));
   mux2X1__0_167 genblk1_17_m8 (.in0(z3[9]), .in1(z3[17]), .sel(shft[3]), 
      .out(z4[17]));
   mux2X1__0_169 genblk1_18_m8 (.in0(z3[10]), .in1(z3[18]), .sel(shft[3]), 
      .out(z4[18]));
   mux2X1__0_171 genblk1_19_m8 (.in0(z3[11]), .in1(z3[19]), .sel(shft[3]), 
      .out(z4[19]));
   mux2X1__0_173 genblk1_20_m8 (.in0(z3[12]), .in1(z3[20]), .sel(shft[3]), 
      .out(z4[20]));
   mux2X1__0_175 genblk1_21_m8 (.in0(z3[13]), .in1(z3[21]), .sel(shft[3]), 
      .out(z4[21]));
   mux2X1__0_177 genblk1_22_m8 (.in0(z3[14]), .in1(z3[22]), .sel(shft[3]), 
      .out(z4[22]));
   mux2X1__0_179 genblk1_23_m8 (.in0(z3[15]), .in1(z3[23]), .sel(shft[3]), 
      .out(z4[23]));
   mux2X1__0_181 genblk1_24_m8 (.in0(z3[16]), .in1(z3[24]), .sel(shft[3]), 
      .out(z4[24]));
   mux2X1__0_183 genblk1_25_m8 (.in0(z3[17]), .in1(z3[25]), .sel(shft[3]), 
      .out(z4[25]));
   mux2X1__0_185 genblk1_26_m8 (.in0(z3[18]), .in1(z3[26]), .sel(shft[3]), 
      .out(z4[26]));
   mux2X1__0_187 genblk1_27_m8 (.in0(z3[19]), .in1(z3[27]), .sel(shft[3]), 
      .out(z4[27]));
   mux2X1__0_189 genblk1_0_m5 (.in0(), .in1(z2[0]), .sel(shft[2]), .out(z3[0]));
   mux2X1__0_191 genblk1_1_m5 (.in0(), .in1(z2[1]), .sel(shft[2]), .out(z3[1]));
   mux2X1__0_193 genblk1_2_m5 (.in0(), .in1(z2[2]), .sel(shft[2]), .out(z3[2]));
   mux2X1__0_195 genblk1_3_m5 (.in0(), .in1(z2[3]), .sel(shft[2]), .out(z3[3]));
   mux2X1__0_197 genblk1_4_m6 (.in0(z2[0]), .in1(z2[4]), .sel(shft[2]), .out(
      z3[4]));
   mux2X1__0_199 genblk1_5_m6 (.in0(z2[1]), .in1(z2[5]), .sel(shft[2]), .out(
      z3[5]));
   mux2X1__0_201 genblk1_6_m6 (.in0(z2[2]), .in1(z2[6]), .sel(shft[2]), .out(
      z3[6]));
   mux2X1__0_203 genblk1_7_m6 (.in0(z2[3]), .in1(z2[7]), .sel(shft[2]), .out(
      z3[7]));
   mux2X1__0_205 genblk1_8_m6 (.in0(z2[4]), .in1(z2[8]), .sel(shft[2]), .out(
      z3[8]));
   mux2X1__0_207 genblk1_9_m6 (.in0(z2[5]), .in1(z2[9]), .sel(shft[2]), .out(
      z3[9]));
   mux2X1__0_209 genblk1_10_m6 (.in0(z2[6]), .in1(z2[10]), .sel(shft[2]), 
      .out(z3[10]));
   mux2X1__0_211 genblk1_11_m6 (.in0(z2[7]), .in1(z2[11]), .sel(shft[2]), 
      .out(z3[11]));
   mux2X1__0_213 genblk1_12_m6 (.in0(z2[8]), .in1(z2[12]), .sel(shft[2]), 
      .out(z3[12]));
   mux2X1__0_215 genblk1_13_m6 (.in0(z2[9]), .in1(z2[13]), .sel(shft[2]), 
      .out(z3[13]));
   mux2X1__0_217 genblk1_14_m6 (.in0(z2[10]), .in1(z2[14]), .sel(shft[2]), 
      .out(z3[14]));
   mux2X1__0_219 genblk1_15_m6 (.in0(z2[11]), .in1(z2[15]), .sel(shft[2]), 
      .out(z3[15]));
   mux2X1__0_221 genblk1_16_m6 (.in0(z2[12]), .in1(z2[16]), .sel(shft[2]), 
      .out(z3[16]));
   mux2X1__0_223 genblk1_17_m6 (.in0(z2[13]), .in1(z2[17]), .sel(shft[2]), 
      .out(z3[17]));
   mux2X1__0_225 genblk1_18_m6 (.in0(z2[14]), .in1(z2[18]), .sel(shft[2]), 
      .out(z3[18]));
   mux2X1__0_227 genblk1_19_m6 (.in0(z2[15]), .in1(z2[19]), .sel(shft[2]), 
      .out(z3[19]));
   mux2X1__0_229 genblk1_20_m6 (.in0(z2[16]), .in1(z2[20]), .sel(shft[2]), 
      .out(z3[20]));
   mux2X1__0_231 genblk1_21_m6 (.in0(z2[17]), .in1(z2[21]), .sel(shft[2]), 
      .out(z3[21]));
   mux2X1__0_233 genblk1_22_m6 (.in0(z2[18]), .in1(z2[22]), .sel(shft[2]), 
      .out(z3[22]));
   mux2X1__0_235 genblk1_23_m6 (.in0(z2[19]), .in1(z2[23]), .sel(shft[2]), 
      .out(z3[23]));
   mux2X1__0_237 genblk1_24_m6 (.in0(z2[20]), .in1(z2[24]), .sel(shft[2]), 
      .out(z3[24]));
   mux2X1__0_239 genblk1_25_m6 (.in0(z2[21]), .in1(z2[25]), .sel(shft[2]), 
      .out(z3[25]));
   mux2X1__0_241 genblk1_26_m6 (.in0(z2[22]), .in1(z2[26]), .sel(shft[2]), 
      .out(z3[26]));
   mux2X1__0_243 genblk1_27_m6 (.in0(z2[23]), .in1(z2[27]), .sel(shft[2]), 
      .out(z3[27]));
   mux2X1__0_245 genblk1_0_m3 (.in0(), .in1(z1[0]), .sel(shft[1]), .out(z2[0]));
   mux2X1__0_247 genblk1_1_m3 (.in0(), .in1(z1[1]), .sel(shft[1]), .out(z2[1]));
   mux2X1__0_249 genblk1_2_m4 (.in0(z1[0]), .in1(z1[2]), .sel(shft[1]), .out(
      z2[2]));
   mux2X1__0_251 genblk1_3_m4 (.in0(z1[1]), .in1(z1[3]), .sel(shft[1]), .out(
      z2[3]));
   mux2X1__0_253 genblk1_4_m4 (.in0(z1[2]), .in1(z1[4]), .sel(shft[1]), .out(
      z2[4]));
   mux2X1__0_255 genblk1_5_m4 (.in0(z1[3]), .in1(z1[5]), .sel(shft[1]), .out(
      z2[5]));
   mux2X1__0_257 genblk1_6_m4 (.in0(z1[4]), .in1(z1[6]), .sel(shft[1]), .out(
      z2[6]));
   mux2X1__0_259 genblk1_7_m4 (.in0(z1[5]), .in1(z1[7]), .sel(shft[1]), .out(
      z2[7]));
   mux2X1__0_261 genblk1_8_m4 (.in0(z1[6]), .in1(z1[8]), .sel(shft[1]), .out(
      z2[8]));
   mux2X1__0_263 genblk1_9_m4 (.in0(z1[7]), .in1(z1[9]), .sel(shft[1]), .out(
      z2[9]));
   mux2X1__0_265 genblk1_10_m4 (.in0(z1[8]), .in1(z1[10]), .sel(shft[1]), 
      .out(z2[10]));
   mux2X1__0_267 genblk1_11_m4 (.in0(z1[9]), .in1(z1[11]), .sel(shft[1]), 
      .out(z2[11]));
   mux2X1__0_269 genblk1_12_m4 (.in0(z1[10]), .in1(z1[12]), .sel(shft[1]), 
      .out(z2[12]));
   mux2X1__0_271 genblk1_13_m4 (.in0(z1[11]), .in1(z1[13]), .sel(shft[1]), 
      .out(z2[13]));
   mux2X1__0_273 genblk1_14_m4 (.in0(z1[12]), .in1(z1[14]), .sel(shft[1]), 
      .out(z2[14]));
   mux2X1__0_275 genblk1_15_m4 (.in0(z1[13]), .in1(z1[15]), .sel(shft[1]), 
      .out(z2[15]));
   mux2X1__0_277 genblk1_16_m4 (.in0(z1[14]), .in1(z1[16]), .sel(shft[1]), 
      .out(z2[16]));
   mux2X1__0_279 genblk1_17_m4 (.in0(z1[15]), .in1(z1[17]), .sel(shft[1]), 
      .out(z2[17]));
   mux2X1__0_281 genblk1_18_m4 (.in0(z1[16]), .in1(z1[18]), .sel(shft[1]), 
      .out(z2[18]));
   mux2X1__0_283 genblk1_19_m4 (.in0(z1[17]), .in1(z1[19]), .sel(shft[1]), 
      .out(z2[19]));
   mux2X1__0_285 genblk1_20_m4 (.in0(z1[18]), .in1(z1[20]), .sel(shft[1]), 
      .out(z2[20]));
   mux2X1__0_287 genblk1_21_m4 (.in0(z1[19]), .in1(z1[21]), .sel(shft[1]), 
      .out(z2[21]));
   mux2X1__0_289 genblk1_22_m4 (.in0(z1[20]), .in1(z1[22]), .sel(shft[1]), 
      .out(z2[22]));
   mux2X1__0_291 genblk1_23_m4 (.in0(z1[21]), .in1(z1[23]), .sel(shft[1]), 
      .out(z2[23]));
   mux2X1__0_293 genblk1_24_m4 (.in0(z1[22]), .in1(z1[24]), .sel(shft[1]), 
      .out(z2[24]));
   mux2X1__0_295 genblk1_25_m4 (.in0(z1[23]), .in1(z1[25]), .sel(shft[1]), 
      .out(z2[25]));
   mux2X1__0_297 genblk1_26_m4 (.in0(z1[24]), .in1(z1[26]), .sel(shft[1]), 
      .out(z2[26]));
   mux2X1__0_299 genblk1_27_m4 (.in0(z1[25]), .in1(z1[27]), .sel(shft[1]), 
      .out(z2[27]));
   mux2X1__0_301 genblk1_0_m1 (.in0(), .in1(in[0]), .sel(shft[0]), .out(z1[0]));
   mux2X1__0_303 genblk1_1_m2 (.in0(in[0]), .in1(in[1]), .sel(shft[0]), .out(
      z1[1]));
   mux2X1__0_305 genblk1_2_m2 (.in0(in[1]), .in1(in[2]), .sel(shft[0]), .out(
      z1[2]));
   mux2X1__0_307 genblk1_3_m2 (.in0(in[2]), .in1(in[3]), .sel(shft[0]), .out(
      z1[3]));
   mux2X1__0_309 genblk1_4_m2 (.in0(in[3]), .in1(in[4]), .sel(shft[0]), .out(
      z1[4]));
   mux2X1__0_311 genblk1_5_m2 (.in0(in[4]), .in1(in[5]), .sel(shft[0]), .out(
      z1[5]));
   mux2X1__0_313 genblk1_6_m2 (.in0(in[5]), .in1(in[6]), .sel(shft[0]), .out(
      z1[6]));
   mux2X1__0_315 genblk1_7_m2 (.in0(in[6]), .in1(in[7]), .sel(shft[0]), .out(
      z1[7]));
   mux2X1__0_317 genblk1_8_m2 (.in0(in[7]), .in1(in[8]), .sel(shft[0]), .out(
      z1[8]));
   mux2X1__0_319 genblk1_9_m2 (.in0(in[8]), .in1(in[9]), .sel(shft[0]), .out(
      z1[9]));
   mux2X1__0_321 genblk1_10_m2 (.in0(in[9]), .in1(in[10]), .sel(shft[0]), 
      .out(z1[10]));
   mux2X1__0_323 genblk1_11_m2 (.in0(in[10]), .in1(in[11]), .sel(shft[0]), 
      .out(z1[11]));
   mux2X1__0_325 genblk1_12_m2 (.in0(in[11]), .in1(in[12]), .sel(shft[0]), 
      .out(z1[12]));
   mux2X1__0_327 genblk1_13_m2 (.in0(in[12]), .in1(in[13]), .sel(shft[0]), 
      .out(z1[13]));
   mux2X1__0_329 genblk1_14_m2 (.in0(in[13]), .in1(in[14]), .sel(shft[0]), 
      .out(z1[14]));
   mux2X1__0_331 genblk1_15_m2 (.in0(in[14]), .in1(in[15]), .sel(shft[0]), 
      .out(z1[15]));
   mux2X1__0_333 genblk1_16_m2 (.in0(in[15]), .in1(in[16]), .sel(shft[0]), 
      .out(z1[16]));
   mux2X1__0_335 genblk1_17_m2 (.in0(in[16]), .in1(in[17]), .sel(shft[0]), 
      .out(z1[17]));
   mux2X1__0_337 genblk1_18_m2 (.in0(in[17]), .in1(in[18]), .sel(shft[0]), 
      .out(z1[18]));
   mux2X1__0_339 genblk1_19_m2 (.in0(in[18]), .in1(in[19]), .sel(shft[0]), 
      .out(z1[19]));
   mux2X1__0_341 genblk1_20_m2 (.in0(in[19]), .in1(in[20]), .sel(shft[0]), 
      .out(z1[20]));
   mux2X1__0_343 genblk1_21_m2 (.in0(in[20]), .in1(in[21]), .sel(shft[0]), 
      .out(z1[21]));
   mux2X1__0_345 genblk1_22_m2 (.in0(in[21]), .in1(in[22]), .sel(shft[0]), 
      .out(z1[22]));
   mux2X1__0_347 genblk1_23_m2 (.in0(in[22]), .in1(in[23]), .sel(shft[0]), 
      .out(z1[23]));
   mux2X1__0_349 genblk1_24_m2 (.in0(in[23]), .in1(in[24]), .sel(shft[0]), 
      .out(z1[24]));
   mux2X1__0_351 genblk1_25_m2 (.in0(in[24]), .in1(in[25]), .sel(shft[0]), 
      .out(z1[25]));
   mux2X1__0_353 genblk1_26_m2 (.in0(in[25]), .in1(in[26]), .sel(shft[0]), 
      .out(z1[26]));
   mux2X1 genblk1_27_m2 (.in0(in[26]), .in1(in[27]), .sel(shft[0]), .out(z1[27]));
endmodule

module datapath__0_72(p_0, p_1, p_2);
   input p_0;
   input [22:0]p_1;
   output [22:0]p_2;

   HA_X1 i_0 (.A(p_0), .B(p_1[0]), .CO(n_0), .S(p_2[0]));
   HA_X1 i_1 (.A(p_1[1]), .B(n_0), .CO(n_1), .S(p_2[1]));
   HA_X1 i_2 (.A(p_1[2]), .B(n_1), .CO(n_2), .S(p_2[2]));
   HA_X1 i_3 (.A(p_1[3]), .B(n_2), .CO(n_3), .S(p_2[3]));
   HA_X1 i_4 (.A(p_1[4]), .B(n_3), .CO(n_4), .S(p_2[4]));
   HA_X1 i_5 (.A(p_1[5]), .B(n_4), .CO(n_5), .S(p_2[5]));
   HA_X1 i_6 (.A(p_1[6]), .B(n_5), .CO(n_6), .S(p_2[6]));
   HA_X1 i_7 (.A(p_1[7]), .B(n_6), .CO(n_7), .S(p_2[7]));
   HA_X1 i_8 (.A(p_1[8]), .B(n_7), .CO(n_8), .S(p_2[8]));
   HA_X1 i_9 (.A(p_1[9]), .B(n_8), .CO(n_9), .S(p_2[9]));
   HA_X1 i_10 (.A(p_1[10]), .B(n_9), .CO(n_10), .S(p_2[10]));
   HA_X1 i_11 (.A(p_1[11]), .B(n_10), .CO(n_11), .S(p_2[11]));
   HA_X1 i_12 (.A(p_1[12]), .B(n_11), .CO(n_12), .S(p_2[12]));
   HA_X1 i_13 (.A(p_1[13]), .B(n_12), .CO(n_13), .S(p_2[13]));
   HA_X1 i_14 (.A(p_1[14]), .B(n_13), .CO(n_14), .S(p_2[14]));
   HA_X1 i_15 (.A(p_1[15]), .B(n_14), .CO(n_15), .S(p_2[15]));
   HA_X1 i_16 (.A(p_1[16]), .B(n_15), .CO(n_16), .S(p_2[16]));
   HA_X1 i_17 (.A(p_1[17]), .B(n_16), .CO(n_17), .S(p_2[17]));
   HA_X1 i_18 (.A(p_1[18]), .B(n_17), .CO(n_18), .S(p_2[18]));
   HA_X1 i_19 (.A(p_1[19]), .B(n_18), .CO(n_19), .S(p_2[19]));
   HA_X1 i_20 (.A(p_1[20]), .B(n_19), .CO(n_20), .S(p_2[20]));
   HA_X1 i_21 (.A(p_1[21]), .B(n_20), .CO(n_21), .S(p_2[21]));
   XOR2_X1 i_22 (.A(p_1[22]), .B(n_21), .Z(p_2[22]));
endmodule

module round(number, M);
   input [27:0]number;
   output [22:0]M;

   wire n_0_0;

   OR3_X1 i_0_0 (.A1(number[0]), .A2(number[1]), .A3(number[2]), .ZN(n_0_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(number[3]), .ZN(n_0));
   datapath__0_72 i_1 (.p_0(n_0), .p_1({number[26], number[25], number[24], 
      number[23], number[22], number[21], number[20], number[19], number[18], 
      number[17], number[16], number[15], number[14], number[13], number[12], 
      number[11], number[10], number[9], number[8], number[7], number[6], 
      number[5], number[4]}), .p_2(M));
endmodule

module block_norm(ES, Co, MS, M, E);
   input [7:0]ES;
   input Co;
   input [27:0]MS;
   output [22:0]M;
   output [7:0]E;

   wire [4:0]Zcount_aux;
   wire [4:0]shift;
   wire [27:0]number;
   wire [27:0]slct;

   zero_counter zc (.M({n_0, MS[26], MS[25], MS[24], MS[23], MS[22], MS[21], 
      MS[20], MS[19], MS[18], MS[17], MS[16], MS[15], MS[14], MS[13], MS[12], 
      MS[11], MS[10], MS[9], MS[8], MS[7], MS[6], MS[5], MS[4], MS[3], MS[2], 
      MS[1], MS[0]}), .Zcount(Zcount_aux));
   exponent exp (.ES(ES), .Co(Co), .Zcount_aux(Zcount_aux), .shift(shift), 
      .E(E));
   n_shift sh (.shft(shift), .in(MS), .out(number));
   round r (.number({uc_0, slct[26], slct[25], slct[24], slct[23], slct[22], 
      slct[21], slct[20], slct[19], slct[18], slct[17], slct[16], slct[15], 
      slct[14], slct[13], slct[12], slct[11], slct[10], slct[9], slct[8], 
      slct[7], slct[6], slct[5], slct[4], slct[3], slct[2], slct[1], slct[0]}), 
      .M(M));
   MUX2_X1 i_0_0 (.A(number[0]), .B(number[1]), .S(Co), .Z(slct[0]));
   MUX2_X1 i_0_1 (.A(number[1]), .B(number[2]), .S(Co), .Z(slct[1]));
   MUX2_X1 i_0_2 (.A(number[2]), .B(number[3]), .S(Co), .Z(slct[2]));
   MUX2_X1 i_0_3 (.A(number[3]), .B(number[4]), .S(Co), .Z(slct[3]));
   MUX2_X1 i_0_4 (.A(number[4]), .B(number[5]), .S(Co), .Z(slct[4]));
   MUX2_X1 i_0_5 (.A(number[5]), .B(number[6]), .S(Co), .Z(slct[5]));
   MUX2_X1 i_0_6 (.A(number[6]), .B(number[7]), .S(Co), .Z(slct[6]));
   MUX2_X1 i_0_7 (.A(number[7]), .B(number[8]), .S(Co), .Z(slct[7]));
   MUX2_X1 i_0_8 (.A(number[8]), .B(number[9]), .S(Co), .Z(slct[8]));
   MUX2_X1 i_0_9 (.A(number[9]), .B(number[10]), .S(Co), .Z(slct[9]));
   MUX2_X1 i_0_10 (.A(number[10]), .B(number[11]), .S(Co), .Z(slct[10]));
   MUX2_X1 i_0_11 (.A(number[11]), .B(number[12]), .S(Co), .Z(slct[11]));
   MUX2_X1 i_0_12 (.A(number[12]), .B(number[13]), .S(Co), .Z(slct[12]));
   MUX2_X1 i_0_13 (.A(number[13]), .B(number[14]), .S(Co), .Z(slct[13]));
   MUX2_X1 i_0_14 (.A(number[14]), .B(number[15]), .S(Co), .Z(slct[14]));
   MUX2_X1 i_0_15 (.A(number[15]), .B(number[16]), .S(Co), .Z(slct[15]));
   MUX2_X1 i_0_16 (.A(number[16]), .B(number[17]), .S(Co), .Z(slct[16]));
   MUX2_X1 i_0_17 (.A(number[17]), .B(number[18]), .S(Co), .Z(slct[17]));
   MUX2_X1 i_0_18 (.A(number[18]), .B(number[19]), .S(Co), .Z(slct[18]));
   MUX2_X1 i_0_19 (.A(number[19]), .B(number[20]), .S(Co), .Z(slct[19]));
   MUX2_X1 i_0_20 (.A(number[20]), .B(number[21]), .S(Co), .Z(slct[20]));
   MUX2_X1 i_0_21 (.A(number[21]), .B(number[22]), .S(Co), .Z(slct[21]));
   MUX2_X1 i_0_22 (.A(number[22]), .B(number[23]), .S(Co), .Z(slct[22]));
   MUX2_X1 i_0_23 (.A(number[23]), .B(number[24]), .S(Co), .Z(slct[23]));
   MUX2_X1 i_0_24 (.A(number[24]), .B(number[25]), .S(Co), .Z(slct[24]));
   MUX2_X1 i_0_25 (.A(number[25]), .B(number[26]), .S(Co), .Z(slct[25]));
   MUX2_X1 i_0_26 (.A(number[26]), .B(number[27]), .S(Co), .Z(slct[26]));
   OR2_X1 i_0_27 (.A1(MS[27]), .A2(Co), .ZN(n_0));
endmodule

module floating_unit(A, B, A_S, result);
   input [31:0]A;
   input [31:0]B;
   input A_S;
   output [31:0]result;

   wire Enable;
   wire [31:0]S;
   wire [36:0]NB;
   wire [36:0]NA;
   wire [1:0]edata;
   wire [27:0]MBsub;
   wire [27:0]MAsub;
   wire SComp;
   wire [27:0]MBnor;
   wire [27:0]MAnor;
   wire [7:0]Enor;
   wire Compnor;
   wire [27:0]MBout;
   wire [27:0]MAout;
   wire [7:0]Eout;
   wire C;
   wire n_0_0;
   wire CO;
   wire [27:0]MS;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;

   n_case nc (.A(A), .B(B), .S(S), .enable(Enable));
   selector sel (.A({uc_0, A[30], A[29], A[28], A[27], A[26], A[25], A[24], 
      A[23], uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, 
      uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23}), .B({uc_24, B[30], B[29], B[28], B[27], B[26], B[25], B[24], 
      B[23], uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, 
      uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, 
      uc_44, uc_45, uc_46, uc_47}), .edata(edata), .NA({uc_48, uc_49, uc_50, 
      uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, NA[27], uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, 
      uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, 
      uc_80, uc_81, uc_82, uc_83}), .NB({uc_84, uc_85, uc_86, uc_87, uc_88, 
      uc_89, uc_90, uc_91, uc_92, NB[27], uc_93, uc_94, uc_95, uc_96, uc_97, 
      uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, 
      uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, 
      uc_116, uc_117, uc_118, uc_119}));
   n_subn nsbn (.A({uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, uc_126, 
      uc_127, uc_128, NA[27], A[22], A[21], A[20], A[19], A[18], A[17], A[16], 
      A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], 
      A[4], A[3], A[2], A[1], A[0], uc_129, uc_130, uc_131, uc_132}), .B({uc_133, 
      uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, NB[27], 
      B[22], B[21], B[20], B[19], B[18], B[17], B[16], B[15], B[14], B[13], 
      B[12], B[11], B[10], B[9], B[8], B[7], B[6], B[5], B[4], B[3], B[2], B[1], 
      B[0], uc_142, uc_143, uc_144, uc_145}), .Comp(SComp), .SA(), .SB(), .EO(), 
      .MA({MAsub[27], MAsub[26], MAsub[25], MAsub[24], MAsub[23], MAsub[22], 
      MAsub[21], MAsub[20], MAsub[19], MAsub[18], MAsub[17], MAsub[16], 
      MAsub[15], MAsub[14], MAsub[13], MAsub[12], MAsub[11], MAsub[10], MAsub[9], 
      MAsub[8], MAsub[7], MAsub[6], MAsub[5], MAsub[4], uc_146, uc_147, uc_148, 
      uc_149}), .MB({MBsub[27], MBsub[26], MBsub[25], MBsub[24], MBsub[23], 
      MBsub[22], MBsub[21], MBsub[20], MBsub[19], MBsub[18], MBsub[17], 
      MBsub[16], MBsub[15], MBsub[14], MBsub[13], MBsub[12], MBsub[11], 
      MBsub[10], MBsub[9], MBsub[8], MBsub[7], MBsub[6], MBsub[5], MBsub[4], 
      uc_150, uc_151, uc_152, uc_153}));
   n_normal nnrm (.A({uc_154, A[30], A[29], A[28], A[27], A[26], A[25], A[24], 
      A[23], NA[27], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], 
      A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
      A[3], A[2], A[1], A[0], uc_155, uc_156, uc_157, uc_158}), .B({uc_159, 
      B[30], B[29], B[28], B[27], B[26], B[25], B[24], B[23], NB[27], B[22], 
      B[21], B[20], B[19], B[18], B[17], B[16], B[15], B[14], B[13], B[12], 
      B[11], B[10], B[9], B[8], B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0], 
      uc_160, uc_161, uc_162, uc_163}), .edata(edata), .SA(), .SB(), .Comp(
      Compnor), .Enor(Enor), .MA({MAnor[27], MAnor[26], MAnor[25], MAnor[24], 
      MAnor[23], MAnor[22], MAnor[21], MAnor[20], MAnor[19], MAnor[18], 
      MAnor[17], MAnor[16], MAnor[15], MAnor[14], MAnor[13], MAnor[12], 
      MAnor[11], MAnor[10], MAnor[9], MAnor[8], MAnor[7], MAnor[6], MAnor[5], 
      MAnor[4], uc_164, uc_165, uc_166, uc_167}), .MB(MBnor));
   mux_adder mxaddr (.SAsub(), .SBsub(), .SComp(SComp), .Esub({A[30], A[29], 
      A[28], A[27], A[26], A[25], A[24], A[23]}), .MAsub({MAsub[27], MAsub[26], 
      MAsub[25], MAsub[24], MAsub[23], MAsub[22], MAsub[21], MAsub[20], 
      MAsub[19], MAsub[18], MAsub[17], MAsub[16], MAsub[15], MAsub[14], 
      MAsub[13], MAsub[12], MAsub[11], MAsub[10], MAsub[9], MAsub[8], MAsub[7], 
      MAsub[6], MAsub[5], MAsub[4], uc_168, uc_169, uc_170, uc_171}), .MBsub({
      MBsub[27], MBsub[26], MBsub[25], MBsub[24], MBsub[23], MBsub[22], 
      MBsub[21], MBsub[20], MBsub[19], MBsub[18], MBsub[17], MBsub[16], 
      MBsub[15], MBsub[14], MBsub[13], MBsub[12], MBsub[11], MBsub[10], MBsub[9], 
      MBsub[8], MBsub[7], MBsub[6], MBsub[5], MBsub[4], uc_172, uc_173, uc_174, 
      uc_175}), .SAnor(), .SBnor(), .NComp(Compnor), .Enor(Enor), .MAnor({
      MAnor[27], MAnor[26], MAnor[25], MAnor[24], MAnor[23], MAnor[22], 
      MAnor[21], MAnor[20], MAnor[19], MAnor[18], MAnor[17], MAnor[16], 
      MAnor[15], MAnor[14], MAnor[13], MAnor[12], MAnor[11], MAnor[10], MAnor[9], 
      MAnor[8], MAnor[7], MAnor[6], MAnor[5], MAnor[4], uc_176, uc_177, uc_178, 
      uc_179}), .MBnor(MBnor), .edata(edata), .SA(), .SB(), .C(C), .Eout(Eout), 
      .MAout({MAout[27], MAout[26], MAout[25], MAout[24], MAout[23], MAout[22], 
      MAout[21], MAout[20], MAout[19], MAout[18], MAout[17], MAout[16], 
      MAout[15], MAout[14], MAout[13], MAout[12], MAout[11], MAout[10], MAout[9], 
      MAout[8], MAout[7], MAout[6], MAout[5], MAout[4], uc_180, uc_181, uc_182, 
      uc_183}), .MBout(MBout));
   block_adder ba (.SA(A[31]), .SB(B[31]), .Comp(C), .A({MAout[27], MAout[26], 
      MAout[25], MAout[24], MAout[23], MAout[22], MAout[21], MAout[20], 
      MAout[19], MAout[18], MAout[17], MAout[16], MAout[15], MAout[14], 
      MAout[13], MAout[12], MAout[11], MAout[10], MAout[9], MAout[8], MAout[7], 
      MAout[6], MAout[5], MAout[4], uc_184, uc_185, uc_186, uc_187}), .B(MBout), 
      .A_S(A_S), .MS(MS), .CO(CO), .SO(n_0_0));
   block_norm blknrm (.ES(Eout), .Co(CO), .MS(MS), .M({n_0_31, n_0_30, n_0_29, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
      n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
      n_0_10, n_0_9}), .E({n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1}));
   MUX2_X1 i_0_0_0 (.A(S[0]), .B(n_0_9), .S(Enable), .Z(result[0]));
   MUX2_X1 i_0_0_1 (.A(S[1]), .B(n_0_10), .S(Enable), .Z(result[1]));
   MUX2_X1 i_0_0_2 (.A(S[2]), .B(n_0_11), .S(Enable), .Z(result[2]));
   MUX2_X1 i_0_0_3 (.A(S[3]), .B(n_0_12), .S(Enable), .Z(result[3]));
   MUX2_X1 i_0_0_4 (.A(S[4]), .B(n_0_13), .S(Enable), .Z(result[4]));
   MUX2_X1 i_0_0_5 (.A(S[5]), .B(n_0_14), .S(Enable), .Z(result[5]));
   MUX2_X1 i_0_0_6 (.A(S[6]), .B(n_0_15), .S(Enable), .Z(result[6]));
   MUX2_X1 i_0_0_7 (.A(S[7]), .B(n_0_16), .S(Enable), .Z(result[7]));
   MUX2_X1 i_0_0_8 (.A(S[8]), .B(n_0_17), .S(Enable), .Z(result[8]));
   MUX2_X1 i_0_0_9 (.A(S[9]), .B(n_0_18), .S(Enable), .Z(result[9]));
   MUX2_X1 i_0_0_10 (.A(S[10]), .B(n_0_19), .S(Enable), .Z(result[10]));
   MUX2_X1 i_0_0_11 (.A(S[11]), .B(n_0_20), .S(Enable), .Z(result[11]));
   MUX2_X1 i_0_0_12 (.A(S[12]), .B(n_0_21), .S(Enable), .Z(result[12]));
   MUX2_X1 i_0_0_13 (.A(S[13]), .B(n_0_22), .S(Enable), .Z(result[13]));
   MUX2_X1 i_0_0_14 (.A(S[14]), .B(n_0_23), .S(Enable), .Z(result[14]));
   MUX2_X1 i_0_0_15 (.A(S[15]), .B(n_0_24), .S(Enable), .Z(result[15]));
   MUX2_X1 i_0_0_16 (.A(S[16]), .B(n_0_25), .S(Enable), .Z(result[16]));
   MUX2_X1 i_0_0_17 (.A(S[17]), .B(n_0_26), .S(Enable), .Z(result[17]));
   MUX2_X1 i_0_0_18 (.A(S[18]), .B(n_0_27), .S(Enable), .Z(result[18]));
   MUX2_X1 i_0_0_19 (.A(S[19]), .B(n_0_28), .S(Enable), .Z(result[19]));
   MUX2_X1 i_0_0_20 (.A(S[20]), .B(n_0_29), .S(Enable), .Z(result[20]));
   MUX2_X1 i_0_0_21 (.A(S[21]), .B(n_0_30), .S(Enable), .Z(result[21]));
   MUX2_X1 i_0_0_22 (.A(S[22]), .B(n_0_31), .S(Enable), .Z(result[22]));
   MUX2_X1 i_0_0_23 (.A(S[23]), .B(n_0_1), .S(Enable), .Z(result[23]));
   MUX2_X1 i_0_0_24 (.A(S[24]), .B(n_0_2), .S(Enable), .Z(result[24]));
   MUX2_X1 i_0_0_25 (.A(S[25]), .B(n_0_3), .S(Enable), .Z(result[25]));
   MUX2_X1 i_0_0_26 (.A(S[26]), .B(n_0_4), .S(Enable), .Z(result[26]));
   MUX2_X1 i_0_0_27 (.A(S[27]), .B(n_0_5), .S(Enable), .Z(result[27]));
   MUX2_X1 i_0_0_28 (.A(S[28]), .B(n_0_6), .S(Enable), .Z(result[28]));
   MUX2_X1 i_0_0_29 (.A(S[29]), .B(n_0_7), .S(Enable), .Z(result[29]));
   MUX2_X1 i_0_0_30 (.A(S[30]), .B(n_0_8), .S(Enable), .Z(result[30]));
   MUX2_X1 i_0_0_31 (.A(S[31]), .B(n_0_0), .S(Enable), .Z(result[31]));
endmodule
