/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Nov  2 22:17:06 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2390341918 */

module halfAdder__0_11(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_12(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_11 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_19(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_20(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_19 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_27(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_24(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_28(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_27 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_24 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_35(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_32(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_36(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_35 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_32 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_43(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_40(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_44(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_43 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_40 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_51(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_48(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_52(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_51 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_48 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_59(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_56(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_60(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_59 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_56 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_67(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_64(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_68(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_67 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_64 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_75(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_72(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_76(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_75 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_72 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_83(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_80(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_84(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_83 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_80 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_91(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_88(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_92(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_91 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_88 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_99(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_96(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_100(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_99 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_96 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_107(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_104(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_108(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_107 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_104 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_115(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_112(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_116(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_115 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_112 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_123(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_120(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_124(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_123 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_120 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_131(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_128(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_132(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_131 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_128 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_139(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_136(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_140(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_139 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_136 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_147(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_144(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_148(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_147 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_144 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_155(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_152(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_156(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_155 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_152 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_163(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_160(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_164(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_163 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_160 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_171(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_168(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_172(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_171 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_168 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_179(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_176(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_180(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_179 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_176 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_187(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_184(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_188(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_187 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_184 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_195(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_192(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_196(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_195 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_192 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_203(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_200(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_204(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_203 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_200 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_211(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_208(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_212(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_211 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_208 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_219(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_216(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_220(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_219 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_216 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_227(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_224(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_228(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_227 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_224 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_235(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_232(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_236(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_235 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_232 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_243(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_240(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_244(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_243 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_240 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_251(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_248(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_252(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_251 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_248 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_259(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_256(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_260(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_259 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_256 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_264(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   XOR2_X1 i_1_0 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_268(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_264 h2d (.in1(y), .in2(cin), .cout(), .sum(sum));
endmodule

module halfAdder__0_275(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_276(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_275 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_283(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_284(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_283 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_291(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_292(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_291 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_299(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_300(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_299 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_307(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_308(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_307 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_315(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_316(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_315 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_323(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_324(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_323 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_331(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_332(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_331 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_339(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_340(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_339 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_347(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_348(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_347 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_355(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_356(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_355 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_363(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_364(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_363 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_371(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_372(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_371 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_379(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_380(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_379 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_387(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_388(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_387 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_395(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_396(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_395 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_403(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_404(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_403 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_411(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_412(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_411 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_419(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_420(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_419 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_427(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_428(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_427 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_435(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_436(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_435 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_443(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_444(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_443 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_451(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_452(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_451 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_459(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_460(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_459 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_467(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_468(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_467 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_475(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_476(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_475 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_483(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_484(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_483 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_491(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_492(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_491 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_499(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_500(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_499 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_507(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_508(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_507 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_4(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_4 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module carrySaveAdder(in1, in2, sum);
   input [31:0]in1;
   input [31:0]in2;
   output [32:0]sum;

   wire [31:0]coutConnectors;
   wire [30:0]cinConnectors;
   wire [30:0]sumConnectors;

   fullAdder__0_12 genblk1_0_FASum (.cin(), .x(in1[0]), .y(in2[0]), .cout(
      coutConnectors[0]), .sum(sum[0]));
   fullAdder__0_20 genblk1_0_FACarry (.cin(), .x(sumConnectors[0]), .y(
      coutConnectors[0]), .cout(cinConnectors[0]), .sum(sum[1]));
   fullAdder__0_28 genblk1_1_FACarry3 (.cin(cinConnectors[0]), .x(
      sumConnectors[1]), .y(coutConnectors[1]), .cout(cinConnectors[1]), 
      .sum(sum[2]));
   fullAdder__0_36 genblk1_2_FACarry3 (.cin(cinConnectors[1]), .x(
      sumConnectors[2]), .y(coutConnectors[2]), .cout(cinConnectors[2]), 
      .sum(sum[3]));
   fullAdder__0_44 genblk1_3_FACarry3 (.cin(cinConnectors[2]), .x(
      sumConnectors[3]), .y(coutConnectors[3]), .cout(cinConnectors[3]), 
      .sum(sum[4]));
   fullAdder__0_52 genblk1_4_FACarry3 (.cin(cinConnectors[3]), .x(
      sumConnectors[4]), .y(coutConnectors[4]), .cout(cinConnectors[4]), 
      .sum(sum[5]));
   fullAdder__0_60 genblk1_5_FACarry3 (.cin(cinConnectors[4]), .x(
      sumConnectors[5]), .y(coutConnectors[5]), .cout(cinConnectors[5]), 
      .sum(sum[6]));
   fullAdder__0_68 genblk1_6_FACarry3 (.cin(cinConnectors[5]), .x(
      sumConnectors[6]), .y(coutConnectors[6]), .cout(cinConnectors[6]), 
      .sum(sum[7]));
   fullAdder__0_76 genblk1_7_FACarry3 (.cin(cinConnectors[6]), .x(
      sumConnectors[7]), .y(coutConnectors[7]), .cout(cinConnectors[7]), 
      .sum(sum[8]));
   fullAdder__0_84 genblk1_8_FACarry3 (.cin(cinConnectors[7]), .x(
      sumConnectors[8]), .y(coutConnectors[8]), .cout(cinConnectors[8]), 
      .sum(sum[9]));
   fullAdder__0_92 genblk1_9_FACarry3 (.cin(cinConnectors[8]), .x(
      sumConnectors[9]), .y(coutConnectors[9]), .cout(cinConnectors[9]), 
      .sum(sum[10]));
   fullAdder__0_100 genblk1_10_FACarry3 (.cin(cinConnectors[9]), .x(
      sumConnectors[10]), .y(coutConnectors[10]), .cout(cinConnectors[10]), 
      .sum(sum[11]));
   fullAdder__0_108 genblk1_11_FACarry3 (.cin(cinConnectors[10]), .x(
      sumConnectors[11]), .y(coutConnectors[11]), .cout(cinConnectors[11]), 
      .sum(sum[12]));
   fullAdder__0_116 genblk1_12_FACarry3 (.cin(cinConnectors[11]), .x(
      sumConnectors[12]), .y(coutConnectors[12]), .cout(cinConnectors[12]), 
      .sum(sum[13]));
   fullAdder__0_124 genblk1_13_FACarry3 (.cin(cinConnectors[12]), .x(
      sumConnectors[13]), .y(coutConnectors[13]), .cout(cinConnectors[13]), 
      .sum(sum[14]));
   fullAdder__0_132 genblk1_14_FACarry3 (.cin(cinConnectors[13]), .x(
      sumConnectors[14]), .y(coutConnectors[14]), .cout(cinConnectors[14]), 
      .sum(sum[15]));
   fullAdder__0_140 genblk1_15_FACarry3 (.cin(cinConnectors[14]), .x(
      sumConnectors[15]), .y(coutConnectors[15]), .cout(cinConnectors[15]), 
      .sum(sum[16]));
   fullAdder__0_148 genblk1_16_FACarry3 (.cin(cinConnectors[15]), .x(
      sumConnectors[16]), .y(coutConnectors[16]), .cout(cinConnectors[16]), 
      .sum(sum[17]));
   fullAdder__0_156 genblk1_17_FACarry3 (.cin(cinConnectors[16]), .x(
      sumConnectors[17]), .y(coutConnectors[17]), .cout(cinConnectors[17]), 
      .sum(sum[18]));
   fullAdder__0_164 genblk1_18_FACarry3 (.cin(cinConnectors[17]), .x(
      sumConnectors[18]), .y(coutConnectors[18]), .cout(cinConnectors[18]), 
      .sum(sum[19]));
   fullAdder__0_172 genblk1_19_FACarry3 (.cin(cinConnectors[18]), .x(
      sumConnectors[19]), .y(coutConnectors[19]), .cout(cinConnectors[19]), 
      .sum(sum[20]));
   fullAdder__0_180 genblk1_20_FACarry3 (.cin(cinConnectors[19]), .x(
      sumConnectors[20]), .y(coutConnectors[20]), .cout(cinConnectors[20]), 
      .sum(sum[21]));
   fullAdder__0_188 genblk1_21_FACarry3 (.cin(cinConnectors[20]), .x(
      sumConnectors[21]), .y(coutConnectors[21]), .cout(cinConnectors[21]), 
      .sum(sum[22]));
   fullAdder__0_196 genblk1_22_FACarry3 (.cin(cinConnectors[21]), .x(
      sumConnectors[22]), .y(coutConnectors[22]), .cout(cinConnectors[22]), 
      .sum(sum[23]));
   fullAdder__0_204 genblk1_23_FACarry3 (.cin(cinConnectors[22]), .x(
      sumConnectors[23]), .y(coutConnectors[23]), .cout(cinConnectors[23]), 
      .sum(sum[24]));
   fullAdder__0_212 genblk1_24_FACarry3 (.cin(cinConnectors[23]), .x(
      sumConnectors[24]), .y(coutConnectors[24]), .cout(cinConnectors[24]), 
      .sum(sum[25]));
   fullAdder__0_220 genblk1_25_FACarry3 (.cin(cinConnectors[24]), .x(
      sumConnectors[25]), .y(coutConnectors[25]), .cout(cinConnectors[25]), 
      .sum(sum[26]));
   fullAdder__0_228 genblk1_26_FACarry3 (.cin(cinConnectors[25]), .x(
      sumConnectors[26]), .y(coutConnectors[26]), .cout(cinConnectors[26]), 
      .sum(sum[27]));
   fullAdder__0_236 genblk1_27_FACarry3 (.cin(cinConnectors[26]), .x(
      sumConnectors[27]), .y(coutConnectors[27]), .cout(cinConnectors[27]), 
      .sum(sum[28]));
   fullAdder__0_244 genblk1_28_FACarry3 (.cin(cinConnectors[27]), .x(
      sumConnectors[28]), .y(coutConnectors[28]), .cout(cinConnectors[28]), 
      .sum(sum[29]));
   fullAdder__0_252 genblk1_29_FACarry3 (.cin(cinConnectors[28]), .x(
      sumConnectors[29]), .y(coutConnectors[29]), .cout(cinConnectors[29]), 
      .sum(sum[30]));
   fullAdder__0_260 genblk1_30_FACarry3 (.cin(cinConnectors[29]), .x(
      sumConnectors[30]), .y(coutConnectors[30]), .cout(cinConnectors[30]), 
      .sum(sum[31]));
   fullAdder__0_268 genblk1_31_FACarry2 (.cin(cinConnectors[30]), .x(), .y(
      coutConnectors[31]), .cout(), .sum(sum[32]));
   fullAdder__0_276 genblk1_1_FASum (.cin(), .x(in1[1]), .y(in2[1]), .cout(
      coutConnectors[1]), .sum(sumConnectors[0]));
   fullAdder__0_284 genblk1_2_FASum (.cin(), .x(in1[2]), .y(in2[2]), .cout(
      coutConnectors[2]), .sum(sumConnectors[1]));
   fullAdder__0_292 genblk1_3_FASum (.cin(), .x(in1[3]), .y(in2[3]), .cout(
      coutConnectors[3]), .sum(sumConnectors[2]));
   fullAdder__0_300 genblk1_4_FASum (.cin(), .x(in1[4]), .y(in2[4]), .cout(
      coutConnectors[4]), .sum(sumConnectors[3]));
   fullAdder__0_308 genblk1_5_FASum (.cin(), .x(in1[5]), .y(in2[5]), .cout(
      coutConnectors[5]), .sum(sumConnectors[4]));
   fullAdder__0_316 genblk1_6_FASum (.cin(), .x(in1[6]), .y(in2[6]), .cout(
      coutConnectors[6]), .sum(sumConnectors[5]));
   fullAdder__0_324 genblk1_7_FASum (.cin(), .x(in1[7]), .y(in2[7]), .cout(
      coutConnectors[7]), .sum(sumConnectors[6]));
   fullAdder__0_332 genblk1_8_FASum (.cin(), .x(in1[8]), .y(in2[8]), .cout(
      coutConnectors[8]), .sum(sumConnectors[7]));
   fullAdder__0_340 genblk1_9_FASum (.cin(), .x(in1[9]), .y(in2[9]), .cout(
      coutConnectors[9]), .sum(sumConnectors[8]));
   fullAdder__0_348 genblk1_10_FASum (.cin(), .x(in1[10]), .y(in2[10]), .cout(
      coutConnectors[10]), .sum(sumConnectors[9]));
   fullAdder__0_356 genblk1_11_FASum (.cin(), .x(in1[11]), .y(in2[11]), .cout(
      coutConnectors[11]), .sum(sumConnectors[10]));
   fullAdder__0_364 genblk1_12_FASum (.cin(), .x(in1[12]), .y(in2[12]), .cout(
      1'b0), .sum(sumConnectors[11]));
   fullAdder__0_372 genblk1_13_FASum (.cin(), .x(in1[13]), .y(in2[13]), .cout(
      1'b0), .sum(sumConnectors[12]));
   fullAdder__0_380 genblk1_14_FASum (.cin(), .x(in1[14]), .y(in2[14]), .cout(
      coutConnectors[14]), .sum(sumConnectors[13]));
   fullAdder__0_388 genblk1_15_FASum (.cin(), .x(in1[15]), .y(in2[15]), .cout(
      coutConnectors[15]), .sum(sumConnectors[14]));
   fullAdder__0_396 genblk1_16_FASum (.cin(), .x(in1[16]), .y(in2[16]), .cout(
      coutConnectors[16]), .sum(sumConnectors[15]));
   fullAdder__0_404 genblk1_17_FASum (.cin(), .x(in1[17]), .y(in2[17]), .cout(
      coutConnectors[17]), .sum(sumConnectors[16]));
   fullAdder__0_412 genblk1_18_FASum (.cin(), .x(in1[18]), .y(in2[18]), .cout(
      coutConnectors[18]), .sum(sumConnectors[17]));
   fullAdder__0_420 genblk1_19_FASum (.cin(), .x(in1[19]), .y(in2[19]), .cout(
      coutConnectors[19]), .sum(sumConnectors[18]));
   fullAdder__0_428 genblk1_20_FASum (.cin(), .x(in1[20]), .y(in2[20]), .cout(
      coutConnectors[20]), .sum(sumConnectors[19]));
   fullAdder__0_436 genblk1_21_FASum (.cin(), .x(in1[21]), .y(in2[21]), .cout(
      coutConnectors[21]), .sum(sumConnectors[20]));
   fullAdder__0_444 genblk1_22_FASum (.cin(), .x(in1[22]), .y(in2[22]), .cout(
      coutConnectors[22]), .sum(sumConnectors[21]));
   fullAdder__0_452 genblk1_23_FASum (.cin(), .x(in1[23]), .y(in2[23]), .cout(
      coutConnectors[23]), .sum(sumConnectors[22]));
   fullAdder__0_460 genblk1_24_FASum (.cin(), .x(in1[24]), .y(in2[24]), .cout(
      coutConnectors[24]), .sum(sumConnectors[23]));
   fullAdder__0_468 genblk1_25_FASum (.cin(), .x(in1[25]), .y(in2[25]), .cout(
      coutConnectors[25]), .sum(sumConnectors[24]));
   fullAdder__0_476 genblk1_26_FASum (.cin(), .x(in1[26]), .y(in2[26]), .cout(
      coutConnectors[26]), .sum(sumConnectors[25]));
   fullAdder__0_484 genblk1_27_FASum (.cin(), .x(in1[27]), .y(in2[27]), .cout(
      coutConnectors[27]), .sum(sumConnectors[26]));
   fullAdder__0_492 genblk1_28_FASum (.cin(), .x(in1[28]), .y(in2[28]), .cout(
      coutConnectors[28]), .sum(sumConnectors[27]));
   fullAdder__0_500 genblk1_29_FASum (.cin(), .x(in1[29]), .y(in2[29]), .cout(
      coutConnectors[29]), .sum(sumConnectors[28]));
   fullAdder__0_508 genblk1_30_FASum (.cin(), .x(in1[30]), .y(in2[30]), .cout(
      coutConnectors[30]), .sum(sumConnectors[29]));
   fullAdder genblk1_31_FASum (.cin(), .x(in1[31]), .y(in2[31]), .cout(
      coutConnectors[31]), .sum(sumConnectors[30]));
endmodule
