/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 17 18:59:25 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2790001319 */

/* blackbox module registerNbits_bbox_0 */

/* blackbox module registerNbits_bbox_1 */

/* blackbox module registerNbits_bbox */

module datapath(p_0, multiplicand);
   output [31:0]p_0;
   input [31:0]multiplicand;

   INV_X1 i_0 (.A(multiplicand[0]), .ZN(n_0));
   XNOR2_X1 i_1 (.A(multiplicand[1]), .B(n_0), .ZN(p_0[1]));
   NOR2_X1 i_2 (.A1(multiplicand[1]), .A2(multiplicand[0]), .ZN(n_1));
   XNOR2_X1 i_3 (.A(multiplicand[2]), .B(n_1), .ZN(p_0[2]));
   NOR2_X1 i_4 (.A1(multiplicand[2]), .A2(n_3), .ZN(n_2));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   XNOR2_X1 i_6 (.A(multiplicand[3]), .B(n_2), .ZN(p_0[3]));
   NOR2_X1 i_7 (.A1(multiplicand[3]), .A2(n_5), .ZN(n_4));
   INV_X1 i_8 (.A(n_2), .ZN(n_5));
   XNOR2_X1 i_9 (.A(multiplicand[4]), .B(n_4), .ZN(p_0[4]));
   NOR2_X1 i_10 (.A1(multiplicand[4]), .A2(n_7), .ZN(n_6));
   INV_X1 i_11 (.A(n_4), .ZN(n_7));
   XNOR2_X1 i_12 (.A(multiplicand[5]), .B(n_6), .ZN(p_0[5]));
   NOR2_X1 i_13 (.A1(multiplicand[5]), .A2(n_9), .ZN(n_8));
   INV_X1 i_14 (.A(n_6), .ZN(n_9));
   XNOR2_X1 i_15 (.A(multiplicand[6]), .B(n_8), .ZN(p_0[6]));
   NOR2_X1 i_16 (.A1(multiplicand[6]), .A2(n_11), .ZN(n_10));
   INV_X1 i_17 (.A(n_8), .ZN(n_11));
   XNOR2_X1 i_18 (.A(multiplicand[7]), .B(n_10), .ZN(p_0[7]));
   NOR2_X1 i_19 (.A1(multiplicand[7]), .A2(n_13), .ZN(n_12));
   INV_X1 i_20 (.A(n_10), .ZN(n_13));
   XNOR2_X1 i_21 (.A(multiplicand[8]), .B(n_12), .ZN(p_0[8]));
   NOR2_X1 i_22 (.A1(multiplicand[8]), .A2(n_15), .ZN(n_14));
   INV_X1 i_23 (.A(n_12), .ZN(n_15));
   XNOR2_X1 i_24 (.A(multiplicand[9]), .B(n_14), .ZN(p_0[9]));
   NOR2_X1 i_25 (.A1(multiplicand[9]), .A2(n_17), .ZN(n_16));
   INV_X1 i_26 (.A(n_14), .ZN(n_17));
   XNOR2_X1 i_27 (.A(multiplicand[10]), .B(n_16), .ZN(p_0[10]));
   NOR2_X1 i_28 (.A1(multiplicand[10]), .A2(n_19), .ZN(n_18));
   INV_X1 i_29 (.A(n_16), .ZN(n_19));
   XNOR2_X1 i_30 (.A(multiplicand[11]), .B(n_18), .ZN(p_0[11]));
   NOR2_X1 i_31 (.A1(multiplicand[11]), .A2(n_21), .ZN(n_20));
   INV_X1 i_32 (.A(n_18), .ZN(n_21));
   XNOR2_X1 i_33 (.A(multiplicand[12]), .B(n_20), .ZN(p_0[12]));
   NOR2_X1 i_34 (.A1(multiplicand[12]), .A2(n_23), .ZN(n_22));
   INV_X1 i_35 (.A(n_20), .ZN(n_23));
   XNOR2_X1 i_36 (.A(multiplicand[13]), .B(n_22), .ZN(p_0[13]));
   NOR2_X1 i_37 (.A1(multiplicand[13]), .A2(n_25), .ZN(n_24));
   INV_X1 i_38 (.A(n_22), .ZN(n_25));
   XNOR2_X1 i_39 (.A(multiplicand[14]), .B(n_24), .ZN(p_0[14]));
   NOR2_X1 i_40 (.A1(multiplicand[14]), .A2(n_27), .ZN(n_26));
   INV_X1 i_41 (.A(n_24), .ZN(n_27));
   XNOR2_X1 i_42 (.A(multiplicand[15]), .B(n_26), .ZN(p_0[15]));
   NOR2_X1 i_43 (.A1(multiplicand[15]), .A2(n_29), .ZN(n_28));
   INV_X1 i_44 (.A(n_26), .ZN(n_29));
   XNOR2_X1 i_45 (.A(multiplicand[16]), .B(n_28), .ZN(p_0[16]));
   NOR2_X1 i_46 (.A1(multiplicand[16]), .A2(n_31), .ZN(n_30));
   INV_X1 i_47 (.A(n_28), .ZN(n_31));
   XNOR2_X1 i_48 (.A(multiplicand[17]), .B(n_30), .ZN(p_0[17]));
   NOR2_X1 i_49 (.A1(multiplicand[17]), .A2(n_33), .ZN(n_32));
   INV_X1 i_50 (.A(n_30), .ZN(n_33));
   XNOR2_X1 i_51 (.A(multiplicand[18]), .B(n_32), .ZN(p_0[18]));
   NOR2_X1 i_52 (.A1(multiplicand[18]), .A2(n_35), .ZN(n_34));
   INV_X1 i_53 (.A(n_32), .ZN(n_35));
   XNOR2_X1 i_54 (.A(multiplicand[19]), .B(n_34), .ZN(p_0[19]));
   NOR2_X1 i_55 (.A1(multiplicand[19]), .A2(n_37), .ZN(n_36));
   INV_X1 i_56 (.A(n_34), .ZN(n_37));
   XNOR2_X1 i_57 (.A(multiplicand[20]), .B(n_36), .ZN(p_0[20]));
   NOR2_X1 i_58 (.A1(multiplicand[20]), .A2(n_39), .ZN(n_38));
   INV_X1 i_59 (.A(n_36), .ZN(n_39));
   XNOR2_X1 i_60 (.A(multiplicand[21]), .B(n_38), .ZN(p_0[21]));
   NOR2_X1 i_61 (.A1(multiplicand[21]), .A2(n_41), .ZN(n_40));
   INV_X1 i_62 (.A(n_38), .ZN(n_41));
   XNOR2_X1 i_63 (.A(multiplicand[22]), .B(n_40), .ZN(p_0[22]));
   NOR2_X1 i_64 (.A1(multiplicand[22]), .A2(n_43), .ZN(n_42));
   INV_X1 i_65 (.A(n_40), .ZN(n_43));
   XNOR2_X1 i_66 (.A(multiplicand[23]), .B(n_42), .ZN(p_0[23]));
   NOR2_X1 i_67 (.A1(multiplicand[23]), .A2(n_45), .ZN(n_44));
   INV_X1 i_68 (.A(n_42), .ZN(n_45));
   XNOR2_X1 i_69 (.A(multiplicand[24]), .B(n_44), .ZN(p_0[24]));
   NOR2_X1 i_70 (.A1(multiplicand[24]), .A2(n_47), .ZN(n_46));
   INV_X1 i_71 (.A(n_44), .ZN(n_47));
   XNOR2_X1 i_72 (.A(multiplicand[25]), .B(n_46), .ZN(p_0[25]));
   NOR2_X1 i_73 (.A1(multiplicand[25]), .A2(n_49), .ZN(n_48));
   INV_X1 i_74 (.A(n_46), .ZN(n_49));
   XNOR2_X1 i_75 (.A(multiplicand[26]), .B(n_48), .ZN(p_0[26]));
   NOR2_X1 i_76 (.A1(multiplicand[26]), .A2(n_51), .ZN(n_50));
   INV_X1 i_77 (.A(n_48), .ZN(n_51));
   XNOR2_X1 i_78 (.A(multiplicand[27]), .B(n_50), .ZN(p_0[27]));
   NOR2_X1 i_79 (.A1(multiplicand[27]), .A2(n_53), .ZN(n_52));
   INV_X1 i_80 (.A(n_50), .ZN(n_53));
   XNOR2_X1 i_81 (.A(multiplicand[28]), .B(n_52), .ZN(p_0[28]));
   NOR2_X1 i_82 (.A1(multiplicand[28]), .A2(n_55), .ZN(n_54));
   INV_X1 i_83 (.A(n_52), .ZN(n_55));
   XNOR2_X1 i_84 (.A(multiplicand[29]), .B(n_54), .ZN(p_0[29]));
   NOR2_X1 i_85 (.A1(multiplicand[29]), .A2(n_57), .ZN(n_56));
   INV_X1 i_86 (.A(n_54), .ZN(n_57));
   XNOR2_X1 i_87 (.A(multiplicand[30]), .B(n_56), .ZN(p_0[30]));
   NOR2_X1 i_88 (.A1(multiplicand[30]), .A2(n_59), .ZN(n_58));
   INV_X1 i_89 (.A(n_56), .ZN(n_59));
   XNOR2_X1 i_90 (.A(multiplicand[31]), .B(n_58), .ZN(p_0[31]));
endmodule

module datapath__0_109(subRes, subRes0, subRes1, subRes2, subRes3, subRes4, 
      subRes5, subRes6, subRes7, subRes8, subRes9, subRes10, subRes11, subRes12, 
      subRes13, subRes14, product_reg);
   input [63:0]subRes;
   input [63:0]subRes0;
   input [63:0]subRes1;
   input [63:0]subRes2;
   input [63:0]subRes3;
   input [63:0]subRes4;
   input [63:0]subRes5;
   input [63:0]subRes6;
   input [63:0]subRes7;
   input [63:0]subRes8;
   input [63:0]subRes9;
   input [63:0]subRes10;
   input [63:0]subRes11;
   input [63:0]subRes12;
   input [63:0]subRes13;
   input [63:0]subRes14;
   output [63:0]product_reg;

   HA_X1 i_0 (.A(subRes[4]), .B(subRes0[4]), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(subRes[5]), .B(subRes0[5]), .CI(subRes14[5]), .CO(n_3), 
      .S(n_2));
   FA_X1 i_2 (.A(subRes[6]), .B(subRes0[6]), .CI(subRes1[6]), .CO(n_5), .S(n_4));
   HA_X1 i_3 (.A(subRes14[6]), .B(n_3), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(subRes[7]), .B(subRes0[7]), .CI(subRes1[7]), .CO(n_9), .S(n_8));
   FA_X1 i_5 (.A(subRes14[7]), .B(n_5), .CI(n_7), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(subRes[8]), .B(subRes0[8]), .CI(subRes1[8]), .CO(n_13), 
      .S(n_12));
   FA_X1 i_7 (.A(subRes2[8]), .B(subRes14[8]), .CI(n_9), .CO(n_15), .S(n_14));
   HA_X1 i_8 (.A(n_11), .B(n_14), .CO(n_17), .S(n_16));
   FA_X1 i_9 (.A(subRes[9]), .B(subRes0[9]), .CI(subRes1[9]), .CO(n_19), 
      .S(n_18));
   FA_X1 i_10 (.A(subRes2[9]), .B(subRes14[9]), .CI(n_13), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(n_15), .B(n_20), .CI(n_18), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(subRes[10]), .B(subRes0[10]), .CI(subRes1[10]), .CO(n_25), 
      .S(n_24));
   FA_X1 i_13 (.A(subRes2[10]), .B(subRes3[10]), .CI(subRes14[10]), .CO(n_27), 
      .S(n_26));
   FA_X1 i_14 (.A(n_19), .B(n_21), .CI(n_26), .CO(n_29), .S(n_28));
   HA_X1 i_15 (.A(n_24), .B(n_23), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(subRes[11]), .B(subRes0[11]), .CI(subRes1[11]), .CO(n_33), 
      .S(n_32));
   FA_X1 i_17 (.A(subRes2[11]), .B(subRes3[11]), .CI(subRes14[11]), .CO(n_35), 
      .S(n_34));
   FA_X1 i_18 (.A(n_27), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_29), .CI(n_36), .CO(n_39), .S(n_38));
   FA_X1 i_20 (.A(subRes[12]), .B(subRes0[12]), .CI(subRes1[12]), .CO(n_41), 
      .S(n_40));
   FA_X1 i_21 (.A(subRes2[12]), .B(subRes3[12]), .CI(subRes4[12]), .CO(n_43), 
      .S(n_42));
   FA_X1 i_22 (.A(subRes14[12]), .B(n_35), .CI(n_33), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(n_42), .B(n_40), .CI(n_44), .CO(n_47), .S(n_46));
   HA_X1 i_24 (.A(n_37), .B(n_39), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(subRes[13]), .B(subRes0[13]), .CI(subRes1[13]), .CO(n_51), 
      .S(n_50));
   FA_X1 i_26 (.A(subRes2[13]), .B(subRes3[13]), .CI(subRes4[13]), .CO(n_53), 
      .S(n_52));
   FA_X1 i_27 (.A(subRes14[13]), .B(n_43), .CI(n_41), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(n_45), .B(n_52), .CI(n_50), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(n_54), .B(n_47), .CI(n_56), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(subRes[14]), .B(subRes0[14]), .CI(subRes1[14]), .CO(n_61), 
      .S(n_60));
   FA_X1 i_31 (.A(subRes2[14]), .B(subRes3[14]), .CI(subRes4[14]), .CO(n_63), 
      .S(n_62));
   FA_X1 i_32 (.A(subRes5[14]), .B(subRes14[14]), .CI(n_53), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_51), .B(n_55), .CI(n_64), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_62), .B(n_60), .CI(n_57), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_66), .B(n_68), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(subRes[15]), .B(subRes0[15]), .CI(subRes1[15]), .CO(n_73), 
      .S(n_72));
   FA_X1 i_37 (.A(subRes2[15]), .B(subRes3[15]), .CI(subRes4[15]), .CO(n_75), 
      .S(n_74));
   FA_X1 i_38 (.A(subRes5[15]), .B(subRes14[15]), .CI(n_63), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(n_61), .B(n_65), .CI(n_76), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_74), .B(n_72), .CI(n_67), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_69), .CI(n_80), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(subRes[16]), .B(subRes0[16]), .CI(subRes1[16]), .CO(n_85), 
      .S(n_84));
   FA_X1 i_43 (.A(subRes2[16]), .B(subRes3[16]), .CI(subRes4[16]), .CO(n_87), 
      .S(n_86));
   FA_X1 i_44 (.A(subRes5[16]), .B(subRes6[16]), .CI(subRes14[16]), .CO(n_89), 
      .S(n_88));
   FA_X1 i_45 (.A(n_75), .B(n_73), .CI(n_77), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(n_88), .B(n_86), .CI(n_84), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(n_90), .B(n_79), .CI(n_81), .CO(n_95), .S(n_94));
   HA_X1 i_48 (.A(n_92), .B(n_94), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(subRes[17]), .B(subRes0[17]), .CI(subRes1[17]), .CO(n_99), 
      .S(n_98));
   FA_X1 i_50 (.A(subRes2[17]), .B(subRes3[17]), .CI(subRes4[17]), .CO(n_101), 
      .S(n_100));
   FA_X1 i_51 (.A(subRes5[17]), .B(subRes6[17]), .CI(subRes14[17]), .CO(n_103), 
      .S(n_102));
   FA_X1 i_52 (.A(n_89), .B(n_87), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_98), .CO(n_107), .S(n_106));
   FA_X1 i_54 (.A(n_91), .B(n_104), .CI(n_93), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(n_106), .B(n_95), .CI(n_108), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(subRes[18]), .B(subRes0[18]), .CI(subRes1[18]), .CO(n_113), 
      .S(n_112));
   FA_X1 i_57 (.A(subRes2[18]), .B(subRes3[18]), .CI(subRes4[18]), .CO(n_115), 
      .S(n_114));
   FA_X1 i_58 (.A(subRes5[18]), .B(subRes6[18]), .CI(subRes7[18]), .CO(n_117), 
      .S(n_116));
   FA_X1 i_59 (.A(subRes14[18]), .B(n_103), .CI(n_101), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_99), .B(n_105), .CI(n_116), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_114), .B(n_112), .CI(n_118), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_107), .B(n_120), .CI(n_109), .CO(n_125), .S(n_124));
   HA_X1 i_63 (.A(n_122), .B(n_124), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(subRes[19]), .B(subRes0[19]), .CI(subRes1[19]), .CO(n_129), 
      .S(n_128));
   FA_X1 i_65 (.A(subRes2[19]), .B(subRes3[19]), .CI(subRes4[19]), .CO(n_131), 
      .S(n_130));
   FA_X1 i_66 (.A(subRes5[19]), .B(subRes6[19]), .CI(subRes7[19]), .CO(n_133), 
      .S(n_132));
   FA_X1 i_67 (.A(subRes14[19]), .B(n_117), .CI(n_115), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(n_113), .B(n_119), .CI(n_132), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(n_130), .B(n_128), .CI(n_134), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(n_121), .B(n_136), .CI(n_123), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_138), .B(n_125), .CI(n_140), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(subRes[20]), .B(subRes0[20]), .CI(subRes1[20]), .CO(n_145), 
      .S(n_144));
   FA_X1 i_73 (.A(subRes2[20]), .B(subRes3[20]), .CI(subRes4[20]), .CO(n_147), 
      .S(n_146));
   FA_X1 i_74 (.A(subRes5[20]), .B(subRes6[20]), .CI(subRes7[20]), .CO(n_149), 
      .S(n_148));
   FA_X1 i_75 (.A(subRes8[20]), .B(subRes14[20]), .CI(n_133), .CO(n_151), 
      .S(n_150));
   FA_X1 i_76 (.A(n_131), .B(n_129), .CI(n_135), .CO(n_153), .S(n_152));
   FA_X1 i_77 (.A(n_150), .B(n_148), .CI(n_146), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(n_144), .B(n_152), .CI(n_137), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(n_139), .B(n_154), .CI(n_141), .CO(n_159), .S(n_158));
   HA_X1 i_80 (.A(n_156), .B(n_158), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(subRes[21]), .B(subRes0[21]), .CI(subRes1[21]), .CO(n_163), 
      .S(n_162));
   FA_X1 i_82 (.A(subRes2[21]), .B(subRes3[21]), .CI(subRes4[21]), .CO(n_165), 
      .S(n_164));
   FA_X1 i_83 (.A(subRes5[21]), .B(subRes6[21]), .CI(subRes7[21]), .CO(n_167), 
      .S(n_166));
   FA_X1 i_84 (.A(subRes8[21]), .B(subRes14[21]), .CI(n_149), .CO(n_169), 
      .S(n_168));
   FA_X1 i_85 (.A(n_147), .B(n_145), .CI(n_151), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_168), .B(n_166), .CI(n_164), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_162), .B(n_153), .CI(n_170), .CO(n_175), .S(n_174));
   FA_X1 i_88 (.A(n_155), .B(n_157), .CI(n_172), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_174), .B(n_159), .CI(n_176), .CO(n_179), .S(n_178));
   FA_X1 i_90 (.A(subRes[22]), .B(subRes0[22]), .CI(subRes1[22]), .CO(n_181), 
      .S(n_180));
   FA_X1 i_91 (.A(subRes2[22]), .B(subRes3[22]), .CI(subRes4[22]), .CO(n_183), 
      .S(n_182));
   FA_X1 i_92 (.A(subRes5[22]), .B(subRes6[22]), .CI(subRes7[22]), .CO(n_185), 
      .S(n_184));
   FA_X1 i_93 (.A(subRes8[22]), .B(subRes9[22]), .CI(subRes14[22]), .CO(n_187), 
      .S(n_186));
   FA_X1 i_94 (.A(n_167), .B(n_165), .CI(n_163), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(n_169), .B(n_186), .CI(n_184), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(n_182), .B(n_180), .CI(n_171), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_188), .B(n_173), .CI(n_175), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_192), .B(n_190), .CI(n_194), .CO(n_197), .S(n_196));
   HA_X1 i_99 (.A(n_177), .B(n_196), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(subRes[23]), .B(subRes0[23]), .CI(subRes1[23]), .CO(n_201), 
      .S(n_200));
   FA_X1 i_101 (.A(subRes2[23]), .B(subRes3[23]), .CI(subRes4[23]), .CO(n_203), 
      .S(n_202));
   FA_X1 i_102 (.A(subRes5[23]), .B(subRes6[23]), .CI(subRes7[23]), .CO(n_205), 
      .S(n_204));
   FA_X1 i_103 (.A(subRes8[23]), .B(subRes9[23]), .CI(subRes14[23]), .CO(n_207), 
      .S(n_206));
   FA_X1 i_104 (.A(n_187), .B(n_185), .CI(n_183), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(n_181), .B(n_189), .CI(n_206), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(n_204), .B(n_202), .CI(n_200), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(n_208), .B(n_191), .CI(n_193), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(n_210), .B(n_212), .CI(n_195), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(n_214), .B(n_197), .CI(n_216), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(subRes[24]), .B(subRes0[24]), .CI(subRes1[24]), .CO(n_221), 
      .S(n_220));
   FA_X1 i_111 (.A(subRes2[24]), .B(subRes3[24]), .CI(subRes4[24]), .CO(n_223), 
      .S(n_222));
   FA_X1 i_112 (.A(subRes5[24]), .B(subRes6[24]), .CI(subRes7[24]), .CO(n_225), 
      .S(n_224));
   FA_X1 i_113 (.A(subRes8[24]), .B(subRes9[24]), .CI(subRes10[24]), .CO(n_227), 
      .S(n_226));
   FA_X1 i_114 (.A(subRes14[24]), .B(n_207), .CI(n_205), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_203), .B(n_201), .CI(n_209), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_226), .B(n_224), .CI(n_222), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_220), .B(n_230), .CI(n_228), .CO(n_235), .S(n_234));
   FA_X1 i_118 (.A(n_213), .B(n_211), .CI(n_215), .CO(n_237), .S(n_236));
   FA_X1 i_119 (.A(n_232), .B(n_236), .CI(n_234), .CO(n_239), .S(n_238));
   HA_X1 i_120 (.A(n_217), .B(n_238), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(subRes[25]), .B(subRes0[25]), .CI(subRes1[25]), .CO(n_243), 
      .S(n_242));
   FA_X1 i_122 (.A(subRes2[25]), .B(subRes3[25]), .CI(subRes4[25]), .CO(n_245), 
      .S(n_244));
   FA_X1 i_123 (.A(subRes5[25]), .B(subRes6[25]), .CI(subRes7[25]), .CO(n_247), 
      .S(n_246));
   FA_X1 i_124 (.A(subRes8[25]), .B(subRes9[25]), .CI(subRes10[25]), .CO(n_249), 
      .S(n_248));
   FA_X1 i_125 (.A(subRes14[25]), .B(n_227), .CI(n_225), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_223), .B(n_221), .CI(n_229), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_248), .B(n_246), .CI(n_244), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_242), .B(n_231), .CI(n_252), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_250), .B(n_233), .CI(n_235), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_254), .B(n_256), .CI(n_237), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_258), .B(n_239), .CI(n_260), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(subRes[26]), .B(subRes0[26]), .CI(subRes1[26]), .CO(n_265), 
      .S(n_264));
   FA_X1 i_133 (.A(subRes2[26]), .B(subRes3[26]), .CI(subRes4[26]), .CO(n_267), 
      .S(n_266));
   FA_X1 i_134 (.A(subRes5[26]), .B(subRes6[26]), .CI(subRes7[26]), .CO(n_269), 
      .S(n_268));
   FA_X1 i_135 (.A(subRes8[26]), .B(subRes9[26]), .CI(subRes10[26]), .CO(n_271), 
      .S(n_270));
   FA_X1 i_136 (.A(subRes11[26]), .B(subRes14[26]), .CI(n_249), .CO(n_273), 
      .S(n_272));
   FA_X1 i_137 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(n_251), .B(n_272), .CI(n_270), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(n_268), .B(n_266), .CI(n_264), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(n_253), .B(n_274), .CI(n_255), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(n_257), .B(n_278), .CI(n_276), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(n_259), .B(n_280), .CI(n_261), .CO(n_285), .S(n_284));
   HA_X1 i_143 (.A(n_282), .B(n_284), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(subRes[27]), .B(subRes0[27]), .CI(subRes1[27]), .CO(n_289), 
      .S(n_288));
   FA_X1 i_145 (.A(subRes2[27]), .B(subRes3[27]), .CI(subRes4[27]), .CO(n_291), 
      .S(n_290));
   FA_X1 i_146 (.A(subRes5[27]), .B(subRes6[27]), .CI(subRes7[27]), .CO(n_293), 
      .S(n_292));
   FA_X1 i_147 (.A(subRes8[27]), .B(subRes9[27]), .CI(subRes10[27]), .CO(n_295), 
      .S(n_294));
   FA_X1 i_148 (.A(subRes11[27]), .B(subRes14[27]), .CI(n_271), .CO(n_297), 
      .S(n_296));
   FA_X1 i_149 (.A(n_269), .B(n_267), .CI(n_265), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_275), .B(n_273), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_294), .B(n_292), .CI(n_290), .CO(n_303), .S(n_302));
   FA_X1 i_152 (.A(n_288), .B(n_298), .CI(n_279), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(n_277), .B(n_300), .CI(n_281), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(n_302), .B(n_304), .CI(n_283), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(n_306), .B(n_285), .CI(n_308), .CO(n_311), .S(n_310));
   FA_X1 i_156 (.A(subRes[28]), .B(subRes0[28]), .CI(subRes1[28]), .CO(n_313), 
      .S(n_312));
   FA_X1 i_157 (.A(subRes2[28]), .B(subRes3[28]), .CI(subRes4[28]), .CO(n_315), 
      .S(n_314));
   FA_X1 i_158 (.A(subRes5[28]), .B(subRes6[28]), .CI(subRes7[28]), .CO(n_317), 
      .S(n_316));
   FA_X1 i_159 (.A(subRes8[28]), .B(subRes9[28]), .CI(subRes10[28]), .CO(n_319), 
      .S(n_318));
   FA_X1 i_160 (.A(subRes11[28]), .B(subRes12[28]), .CI(subRes14[28]), .CO(n_321), 
      .S(n_320));
   FA_X1 i_161 (.A(n_295), .B(n_293), .CI(n_291), .CO(n_323), .S(n_322));
   FA_X1 i_162 (.A(n_289), .B(n_299), .CI(n_297), .CO(n_325), .S(n_324));
   FA_X1 i_163 (.A(n_320), .B(n_318), .CI(n_316), .CO(n_327), .S(n_326));
   FA_X1 i_164 (.A(n_314), .B(n_312), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_165 (.A(n_303), .B(n_301), .CI(n_324), .CO(n_331), .S(n_330));
   FA_X1 i_166 (.A(n_305), .B(n_328), .CI(n_326), .CO(n_333), .S(n_332));
   FA_X1 i_167 (.A(n_307), .B(n_330), .CI(n_309), .CO(n_335), .S(n_334));
   HA_X1 i_168 (.A(n_332), .B(n_334), .CO(n_337), .S(n_336));
   FA_X1 i_169 (.A(subRes[29]), .B(subRes0[29]), .CI(subRes1[29]), .CO(n_339), 
      .S(n_338));
   FA_X1 i_170 (.A(subRes2[29]), .B(subRes3[29]), .CI(subRes4[29]), .CO(n_341), 
      .S(n_340));
   FA_X1 i_171 (.A(subRes5[29]), .B(subRes6[29]), .CI(subRes7[29]), .CO(n_343), 
      .S(n_342));
   FA_X1 i_172 (.A(subRes8[29]), .B(subRes9[29]), .CI(subRes10[29]), .CO(n_345), 
      .S(n_344));
   FA_X1 i_173 (.A(subRes11[29]), .B(subRes12[29]), .CI(subRes14[29]), .CO(n_347), 
      .S(n_346));
   FA_X1 i_174 (.A(n_321), .B(n_319), .CI(n_317), .CO(n_349), .S(n_348));
   FA_X1 i_175 (.A(n_315), .B(n_313), .CI(n_323), .CO(n_351), .S(n_350));
   FA_X1 i_176 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_353), .S(n_352));
   FA_X1 i_177 (.A(n_340), .B(n_338), .CI(n_325), .CO(n_355), .S(n_354));
   FA_X1 i_178 (.A(n_350), .B(n_348), .CI(n_327), .CO(n_357), .S(n_356));
   FA_X1 i_179 (.A(n_329), .B(n_354), .CI(n_352), .CO(n_359), .S(n_358));
   FA_X1 i_180 (.A(n_331), .B(n_356), .CI(n_333), .CO(n_361), .S(n_360));
   FA_X1 i_181 (.A(n_358), .B(n_335), .CI(n_360), .CO(n_363), .S(n_362));
   FA_X1 i_182 (.A(subRes[30]), .B(subRes0[30]), .CI(subRes1[30]), .CO(n_365), 
      .S(n_364));
   FA_X1 i_183 (.A(subRes2[30]), .B(subRes3[30]), .CI(subRes4[30]), .CO(n_367), 
      .S(n_366));
   FA_X1 i_184 (.A(subRes5[30]), .B(subRes6[30]), .CI(subRes7[30]), .CO(n_369), 
      .S(n_368));
   FA_X1 i_185 (.A(subRes8[30]), .B(subRes9[30]), .CI(subRes10[30]), .CO(n_371), 
      .S(n_370));
   FA_X1 i_186 (.A(subRes11[30]), .B(subRes12[30]), .CI(subRes13[30]), .CO(n_373), 
      .S(n_372));
   FA_X1 i_187 (.A(subRes14[30]), .B(n_347), .CI(n_345), .CO(n_375), .S(n_374));
   FA_X1 i_188 (.A(n_343), .B(n_341), .CI(n_339), .CO(n_377), .S(n_376));
   FA_X1 i_189 (.A(n_349), .B(n_372), .CI(n_370), .CO(n_379), .S(n_378));
   FA_X1 i_190 (.A(n_368), .B(n_366), .CI(n_364), .CO(n_381), .S(n_380));
   FA_X1 i_191 (.A(n_351), .B(n_376), .CI(n_374), .CO(n_383), .S(n_382));
   FA_X1 i_192 (.A(n_353), .B(n_355), .CI(n_357), .CO(n_385), .S(n_384));
   FA_X1 i_193 (.A(n_380), .B(n_378), .CI(n_382), .CO(n_387), .S(n_386));
   FA_X1 i_194 (.A(n_359), .B(n_384), .CI(n_361), .CO(n_389), .S(n_388));
   HA_X1 i_195 (.A(n_386), .B(n_388), .CO(n_391), .S(n_390));
   FA_X1 i_196 (.A(subRes[31]), .B(subRes0[31]), .CI(subRes1[31]), .CO(n_393), 
      .S(n_392));
   FA_X1 i_197 (.A(subRes2[31]), .B(subRes3[31]), .CI(subRes4[31]), .CO(n_395), 
      .S(n_394));
   FA_X1 i_198 (.A(subRes5[31]), .B(subRes6[31]), .CI(subRes7[31]), .CO(n_397), 
      .S(n_396));
   FA_X1 i_199 (.A(subRes8[31]), .B(subRes9[31]), .CI(subRes10[31]), .CO(n_399), 
      .S(n_398));
   FA_X1 i_200 (.A(subRes11[31]), .B(subRes12[31]), .CI(subRes13[31]), .CO(n_401), 
      .S(n_400));
   FA_X1 i_201 (.A(subRes14[31]), .B(n_373), .CI(n_371), .CO(n_403), .S(n_402));
   FA_X1 i_202 (.A(n_369), .B(n_367), .CI(n_365), .CO(n_405), .S(n_404));
   FA_X1 i_203 (.A(n_377), .B(n_375), .CI(n_400), .CO(n_407), .S(n_406));
   FA_X1 i_204 (.A(n_398), .B(n_396), .CI(n_394), .CO(n_409), .S(n_408));
   FA_X1 i_205 (.A(n_392), .B(n_404), .CI(n_402), .CO(n_411), .S(n_410));
   FA_X1 i_206 (.A(n_381), .B(n_379), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_207 (.A(n_383), .B(n_408), .CI(n_385), .CO(n_415), .S(n_414));
   FA_X1 i_208 (.A(n_412), .B(n_410), .CI(n_387), .CO(n_417), .S(n_416));
   FA_X1 i_209 (.A(n_414), .B(n_389), .CI(n_416), .CO(n_419), .S(n_418));
   XNOR2_X1 i_210 (.A(subRes[32]), .B(subRes0[32]), .ZN(n_420));
   OR2_X1 i_211 (.A1(subRes[32]), .A2(subRes0[32]), .ZN(n_421));
   FA_X1 i_212 (.A(subRes1[32]), .B(subRes2[32]), .CI(subRes3[32]), .CO(n_423), 
      .S(n_422));
   FA_X1 i_213 (.A(subRes4[32]), .B(subRes5[32]), .CI(subRes6[32]), .CO(n_425), 
      .S(n_424));
   FA_X1 i_214 (.A(subRes7[32]), .B(subRes8[32]), .CI(subRes9[32]), .CO(n_427), 
      .S(n_426));
   FA_X1 i_215 (.A(subRes10[32]), .B(subRes11[32]), .CI(subRes12[32]), .CO(n_429), 
      .S(n_428));
   XNOR2_X1 i_216 (.A(subRes13[32]), .B(subRes14[32]), .ZN(n_430));
   XNOR2_X1 i_217 (.A(n_430), .B(n_401), .ZN(n_431));
   INV_X1 i_218 (.A(n_431), .ZN(n_432));
   NAND3_X1 i_219 (.A1(n_434), .A2(n_436), .A3(n_437), .ZN(n_433));
   NAND2_X1 i_220 (.A1(subRes13[32]), .A2(n_435), .ZN(n_434));
   INV_X1 i_221 (.A(subRes14[32]), .ZN(n_435));
   NAND2_X1 i_222 (.A1(n_401), .A2(subRes13[32]), .ZN(n_436));
   NAND2_X1 i_223 (.A1(n_401), .A2(n_435), .ZN(n_437));
   FA_X1 i_224 (.A(n_399), .B(n_397), .CI(n_395), .CO(n_439), .S(n_438));
   FA_X1 i_225 (.A(n_393), .B(n_405), .CI(n_403), .CO(n_441), .S(n_440));
   FA_X1 i_226 (.A(n_432), .B(n_428), .CI(n_426), .CO(n_443), .S(n_442));
   FA_X1 i_227 (.A(n_424), .B(n_422), .CI(n_420), .CO(n_445), .S(n_444));
   FA_X1 i_228 (.A(n_438), .B(n_409), .CI(n_407), .CO(n_447), .S(n_446));
   FA_X1 i_229 (.A(n_440), .B(n_411), .CI(n_444), .CO(n_449), .S(n_448));
   FA_X1 i_230 (.A(n_442), .B(n_413), .CI(n_446), .CO(n_451), .S(n_450));
   FA_X1 i_231 (.A(n_415), .B(n_448), .CI(n_450), .CO(n_453), .S(n_452));
   HA_X1 i_232 (.A(n_417), .B(n_452), .CO(n_455), .S(n_454));
   XNOR2_X1 i_233 (.A(subRes[33]), .B(subRes0[33]), .ZN(n_456));
   OR2_X1 i_234 (.A1(subRes[33]), .A2(subRes0[33]), .ZN(n_457));
   FA_X1 i_235 (.A(subRes1[33]), .B(subRes2[33]), .CI(subRes3[33]), .CO(n_459), 
      .S(n_458));
   FA_X1 i_236 (.A(subRes4[33]), .B(subRes5[33]), .CI(subRes6[33]), .CO(n_461), 
      .S(n_460));
   FA_X1 i_237 (.A(subRes7[33]), .B(subRes8[33]), .CI(subRes9[33]), .CO(n_463), 
      .S(n_462));
   FA_X1 i_238 (.A(subRes10[33]), .B(subRes11[33]), .CI(subRes12[33]), .CO(n_465), 
      .S(n_464));
   FA_X1 i_239 (.A(subRes13[33]), .B(n_429), .CI(n_427), .CO(n_467), .S(n_466));
   FA_X1 i_240 (.A(n_425), .B(n_423), .CI(n_421), .CO(n_469), .S(n_468));
   FA_X1 i_241 (.A(n_439), .B(n_433), .CI(n_464), .CO(n_471), .S(n_470));
   FA_X1 i_242 (.A(n_462), .B(n_460), .CI(n_458), .CO(n_473), .S(n_472));
   FA_X1 i_243 (.A(n_456), .B(n_441), .CI(n_468), .CO(n_475), .S(n_474));
   FA_X1 i_244 (.A(n_466), .B(n_445), .CI(n_443), .CO(n_477), .S(n_476));
   FA_X1 i_245 (.A(n_470), .B(n_447), .CI(n_472), .CO(n_479), .S(n_478));
   FA_X1 i_246 (.A(n_474), .B(n_476), .CI(n_449), .CO(n_481), .S(n_480));
   FA_X1 i_247 (.A(n_478), .B(n_451), .CI(n_480), .CO(n_483), .S(n_482));
   HA_X1 i_248 (.A(n_453), .B(n_482), .CO(n_485), .S(n_484));
   XNOR2_X1 i_249 (.A(subRes[34]), .B(subRes0[34]), .ZN(n_486));
   XNOR2_X1 i_250 (.A(n_486), .B(subRes1[34]), .ZN(n_487));
   INV_X1 i_251 (.A(n_487), .ZN(n_488));
   NAND3_X1 i_252 (.A1(n_490), .A2(n_492), .A3(n_493), .ZN(n_489));
   NAND2_X1 i_253 (.A1(subRes0[34]), .A2(n_491), .ZN(n_490));
   INV_X1 i_254 (.A(subRes[34]), .ZN(n_491));
   NAND2_X1 i_255 (.A1(subRes1[34]), .A2(n_491), .ZN(n_492));
   NAND2_X1 i_256 (.A1(subRes1[34]), .A2(subRes0[34]), .ZN(n_493));
   FA_X1 i_257 (.A(subRes2[34]), .B(subRes3[34]), .CI(subRes4[34]), .CO(n_495), 
      .S(n_494));
   FA_X1 i_258 (.A(subRes5[34]), .B(subRes6[34]), .CI(subRes7[34]), .CO(n_497), 
      .S(n_496));
   FA_X1 i_259 (.A(subRes8[34]), .B(subRes9[34]), .CI(subRes10[34]), .CO(n_499), 
      .S(n_498));
   FA_X1 i_260 (.A(subRes11[34]), .B(subRes12[34]), .CI(subRes13[34]), .CO(n_501), 
      .S(n_500));
   FA_X1 i_261 (.A(n_465), .B(n_463), .CI(n_461), .CO(n_503), .S(n_502));
   FA_X1 i_262 (.A(n_459), .B(n_457), .CI(n_469), .CO(n_505), .S(n_504));
   FA_X1 i_263 (.A(n_467), .B(n_500), .CI(n_498), .CO(n_507), .S(n_506));
   FA_X1 i_264 (.A(n_496), .B(n_494), .CI(n_488), .CO(n_509), .S(n_508));
   FA_X1 i_265 (.A(n_504), .B(n_502), .CI(n_473), .CO(n_511), .S(n_510));
   FA_X1 i_266 (.A(n_471), .B(n_477), .CI(n_475), .CO(n_513), .S(n_512));
   FA_X1 i_267 (.A(n_508), .B(n_506), .CI(n_510), .CO(n_515), .S(n_514));
   FA_X1 i_268 (.A(n_479), .B(n_512), .CI(n_481), .CO(n_517), .S(n_516));
   FA_X1 i_269 (.A(n_514), .B(n_516), .CI(n_483), .CO(n_519), .S(n_518));
   XNOR2_X1 i_270 (.A(subRes0[35]), .B(subRes1[35]), .ZN(n_520));
   OR2_X1 i_271 (.A1(subRes0[35]), .A2(subRes1[35]), .ZN(n_521));
   FA_X1 i_272 (.A(subRes2[35]), .B(subRes3[35]), .CI(subRes4[35]), .CO(n_523), 
      .S(n_522));
   FA_X1 i_273 (.A(subRes5[35]), .B(subRes6[35]), .CI(subRes7[35]), .CO(n_525), 
      .S(n_524));
   FA_X1 i_274 (.A(subRes8[35]), .B(subRes9[35]), .CI(subRes10[35]), .CO(n_527), 
      .S(n_526));
   FA_X1 i_275 (.A(subRes11[35]), .B(subRes12[35]), .CI(subRes13[35]), .CO(n_529), 
      .S(n_528));
   FA_X1 i_276 (.A(n_501), .B(n_499), .CI(n_497), .CO(n_531), .S(n_530));
   FA_X1 i_277 (.A(n_495), .B(n_489), .CI(n_503), .CO(n_533), .S(n_532));
   FA_X1 i_278 (.A(n_528), .B(n_526), .CI(n_524), .CO(n_535), .S(n_534));
   FA_X1 i_279 (.A(n_522), .B(n_520), .CI(n_505), .CO(n_537), .S(n_536));
   FA_X1 i_280 (.A(n_532), .B(n_530), .CI(n_509), .CO(n_539), .S(n_538));
   FA_X1 i_281 (.A(n_507), .B(n_511), .CI(n_536), .CO(n_541), .S(n_540));
   FA_X1 i_282 (.A(n_534), .B(n_513), .CI(n_538), .CO(n_543), .S(n_542));
   FA_X1 i_283 (.A(n_540), .B(n_515), .CI(n_542), .CO(n_545), .S(n_544));
   HA_X1 i_284 (.A(n_517), .B(n_544), .CO(n_547), .S(n_546));
   XNOR2_X1 i_285 (.A(subRes0[36]), .B(subRes1[36]), .ZN(n_548));
   XNOR2_X1 i_286 (.A(n_548), .B(subRes2[36]), .ZN(n_549));
   INV_X1 i_287 (.A(n_549), .ZN(n_550));
   NAND3_X1 i_288 (.A1(n_552), .A2(n_554), .A3(n_555), .ZN(n_551));
   NAND2_X1 i_289 (.A1(subRes1[36]), .A2(n_553), .ZN(n_552));
   INV_X1 i_290 (.A(subRes0[36]), .ZN(n_553));
   NAND2_X1 i_291 (.A1(subRes2[36]), .A2(n_553), .ZN(n_554));
   NAND2_X1 i_292 (.A1(subRes2[36]), .A2(subRes1[36]), .ZN(n_555));
   FA_X1 i_293 (.A(subRes3[36]), .B(subRes4[36]), .CI(subRes5[36]), .CO(n_557), 
      .S(n_556));
   FA_X1 i_294 (.A(subRes6[36]), .B(subRes7[36]), .CI(subRes8[36]), .CO(n_559), 
      .S(n_558));
   FA_X1 i_295 (.A(subRes9[36]), .B(subRes10[36]), .CI(subRes11[36]), .CO(n_561), 
      .S(n_560));
   FA_X1 i_296 (.A(subRes12[36]), .B(subRes13[36]), .CI(n_529), .CO(n_563), 
      .S(n_562));
   FA_X1 i_297 (.A(n_527), .B(n_525), .CI(n_523), .CO(n_565), .S(n_564));
   FA_X1 i_298 (.A(n_521), .B(n_531), .CI(n_562), .CO(n_567), .S(n_566));
   FA_X1 i_299 (.A(n_560), .B(n_558), .CI(n_556), .CO(n_569), .S(n_568));
   FA_X1 i_300 (.A(n_550), .B(n_533), .CI(n_564), .CO(n_571), .S(n_570));
   FA_X1 i_301 (.A(n_535), .B(n_537), .CI(n_566), .CO(n_573), .S(n_572));
   FA_X1 i_302 (.A(n_539), .B(n_568), .CI(n_570), .CO(n_575), .S(n_574));
   FA_X1 i_303 (.A(n_541), .B(n_572), .CI(n_543), .CO(n_577), .S(n_576));
   FA_X1 i_304 (.A(n_574), .B(n_576), .CI(n_545), .CO(n_579), .S(n_578));
   XNOR2_X1 i_305 (.A(subRes1[37]), .B(subRes2[37]), .ZN(n_580));
   OR2_X1 i_306 (.A1(subRes1[37]), .A2(subRes2[37]), .ZN(n_581));
   FA_X1 i_307 (.A(subRes3[37]), .B(subRes4[37]), .CI(subRes5[37]), .CO(n_583), 
      .S(n_582));
   FA_X1 i_308 (.A(subRes6[37]), .B(subRes7[37]), .CI(subRes8[37]), .CO(n_585), 
      .S(n_584));
   FA_X1 i_309 (.A(subRes9[37]), .B(subRes10[37]), .CI(subRes11[37]), .CO(n_587), 
      .S(n_586));
   FA_X1 i_310 (.A(subRes12[37]), .B(subRes13[37]), .CI(n_561), .CO(n_589), 
      .S(n_588));
   FA_X1 i_311 (.A(n_559), .B(n_557), .CI(n_551), .CO(n_591), .S(n_590));
   FA_X1 i_312 (.A(n_565), .B(n_563), .CI(n_588), .CO(n_593), .S(n_592));
   FA_X1 i_313 (.A(n_586), .B(n_584), .CI(n_582), .CO(n_595), .S(n_594));
   FA_X1 i_314 (.A(n_580), .B(n_590), .CI(n_569), .CO(n_597), .S(n_596));
   FA_X1 i_315 (.A(n_567), .B(n_592), .CI(n_571), .CO(n_599), .S(n_598));
   FA_X1 i_316 (.A(n_594), .B(n_573), .CI(n_596), .CO(n_601), .S(n_600));
   FA_X1 i_317 (.A(n_575), .B(n_598), .CI(n_600), .CO(n_603), .S(n_602));
   HA_X1 i_318 (.A(n_577), .B(n_602), .CO(n_605), .S(n_604));
   XNOR2_X1 i_319 (.A(subRes1[38]), .B(subRes2[38]), .ZN(n_606));
   XNOR2_X1 i_320 (.A(n_606), .B(subRes3[38]), .ZN(n_607));
   INV_X1 i_321 (.A(n_607), .ZN(n_608));
   NAND3_X1 i_322 (.A1(n_610), .A2(n_612), .A3(n_613), .ZN(n_609));
   NAND2_X1 i_323 (.A1(subRes2[38]), .A2(n_611), .ZN(n_610));
   INV_X1 i_324 (.A(subRes1[38]), .ZN(n_611));
   NAND2_X1 i_325 (.A1(subRes3[38]), .A2(n_611), .ZN(n_612));
   NAND2_X1 i_326 (.A1(subRes3[38]), .A2(subRes2[38]), .ZN(n_613));
   FA_X1 i_327 (.A(subRes4[38]), .B(subRes5[38]), .CI(subRes6[38]), .CO(n_615), 
      .S(n_614));
   FA_X1 i_328 (.A(subRes7[38]), .B(subRes8[38]), .CI(subRes9[38]), .CO(n_617), 
      .S(n_616));
   FA_X1 i_329 (.A(subRes10[38]), .B(subRes11[38]), .CI(subRes12[38]), .CO(n_619), 
      .S(n_618));
   FA_X1 i_330 (.A(subRes13[38]), .B(n_587), .CI(n_585), .CO(n_621), .S(n_620));
   FA_X1 i_331 (.A(n_583), .B(n_581), .CI(n_591), .CO(n_623), .S(n_622));
   FA_X1 i_332 (.A(n_589), .B(n_618), .CI(n_616), .CO(n_625), .S(n_624));
   FA_X1 i_333 (.A(n_614), .B(n_608), .CI(n_622), .CO(n_627), .S(n_626));
   FA_X1 i_334 (.A(n_620), .B(n_595), .CI(n_593), .CO(n_629), .S(n_628));
   FA_X1 i_335 (.A(n_597), .B(n_626), .CI(n_624), .CO(n_631), .S(n_630));
   FA_X1 i_336 (.A(n_599), .B(n_628), .CI(n_601), .CO(n_633), .S(n_632));
   FA_X1 i_337 (.A(n_630), .B(n_632), .CI(n_603), .CO(n_635), .S(n_634));
   XNOR2_X1 i_338 (.A(subRes2[39]), .B(subRes3[39]), .ZN(n_636));
   OR2_X1 i_339 (.A1(subRes2[39]), .A2(subRes3[39]), .ZN(n_637));
   FA_X1 i_340 (.A(subRes4[39]), .B(subRes5[39]), .CI(subRes6[39]), .CO(n_639), 
      .S(n_638));
   FA_X1 i_341 (.A(subRes7[39]), .B(subRes8[39]), .CI(subRes9[39]), .CO(n_641), 
      .S(n_640));
   FA_X1 i_342 (.A(subRes10[39]), .B(subRes11[39]), .CI(subRes12[39]), .CO(n_643), 
      .S(n_642));
   FA_X1 i_343 (.A(subRes13[39]), .B(n_619), .CI(n_617), .CO(n_645), .S(n_644));
   FA_X1 i_344 (.A(n_615), .B(n_609), .CI(n_621), .CO(n_647), .S(n_646));
   FA_X1 i_345 (.A(n_642), .B(n_640), .CI(n_638), .CO(n_649), .S(n_648));
   FA_X1 i_346 (.A(n_636), .B(n_623), .CI(n_646), .CO(n_651), .S(n_650));
   FA_X1 i_347 (.A(n_644), .B(n_625), .CI(n_629), .CO(n_653), .S(n_652));
   FA_X1 i_348 (.A(n_627), .B(n_648), .CI(n_650), .CO(n_655), .S(n_654));
   FA_X1 i_349 (.A(n_652), .B(n_631), .CI(n_654), .CO(n_657), .S(n_656));
   HA_X1 i_350 (.A(n_633), .B(n_656), .CO(n_659), .S(n_658));
   XNOR2_X1 i_351 (.A(subRes2[40]), .B(subRes3[40]), .ZN(n_660));
   XNOR2_X1 i_352 (.A(n_660), .B(subRes4[40]), .ZN(n_661));
   INV_X1 i_353 (.A(n_661), .ZN(n_662));
   NAND3_X1 i_354 (.A1(n_664), .A2(n_666), .A3(n_667), .ZN(n_663));
   NAND2_X1 i_355 (.A1(subRes3[40]), .A2(n_665), .ZN(n_664));
   INV_X1 i_356 (.A(subRes2[40]), .ZN(n_665));
   NAND2_X1 i_357 (.A1(subRes4[40]), .A2(n_665), .ZN(n_666));
   NAND2_X1 i_358 (.A1(subRes4[40]), .A2(subRes3[40]), .ZN(n_667));
   FA_X1 i_359 (.A(subRes5[40]), .B(subRes6[40]), .CI(subRes7[40]), .CO(n_669), 
      .S(n_668));
   FA_X1 i_360 (.A(subRes8[40]), .B(subRes9[40]), .CI(subRes10[40]), .CO(n_671), 
      .S(n_670));
   FA_X1 i_361 (.A(subRes11[40]), .B(subRes12[40]), .CI(subRes13[40]), .CO(n_673), 
      .S(n_672));
   FA_X1 i_362 (.A(n_643), .B(n_641), .CI(n_639), .CO(n_675), .S(n_674));
   FA_X1 i_363 (.A(n_637), .B(n_645), .CI(n_672), .CO(n_677), .S(n_676));
   FA_X1 i_364 (.A(n_670), .B(n_668), .CI(n_662), .CO(n_679), .S(n_678));
   FA_X1 i_365 (.A(n_647), .B(n_674), .CI(n_649), .CO(n_681), .S(n_680));
   FA_X1 i_366 (.A(n_676), .B(n_651), .CI(n_678), .CO(n_683), .S(n_682));
   FA_X1 i_367 (.A(n_653), .B(n_680), .CI(n_655), .CO(n_685), .S(n_684));
   FA_X1 i_368 (.A(n_682), .B(n_684), .CI(n_657), .CO(n_687), .S(n_686));
   XNOR2_X1 i_369 (.A(subRes3[41]), .B(subRes4[41]), .ZN(n_688));
   OR2_X1 i_370 (.A1(subRes3[41]), .A2(subRes4[41]), .ZN(n_689));
   FA_X1 i_371 (.A(subRes5[41]), .B(subRes6[41]), .CI(subRes7[41]), .CO(n_691), 
      .S(n_690));
   FA_X1 i_372 (.A(subRes8[41]), .B(subRes9[41]), .CI(subRes10[41]), .CO(n_693), 
      .S(n_692));
   FA_X1 i_373 (.A(subRes11[41]), .B(subRes12[41]), .CI(subRes13[41]), .CO(n_695), 
      .S(n_694));
   FA_X1 i_374 (.A(n_673), .B(n_671), .CI(n_669), .CO(n_697), .S(n_696));
   FA_X1 i_375 (.A(n_663), .B(n_675), .CI(n_694), .CO(n_699), .S(n_698));
   FA_X1 i_376 (.A(n_692), .B(n_690), .CI(n_688), .CO(n_701), .S(n_700));
   FA_X1 i_377 (.A(n_696), .B(n_679), .CI(n_677), .CO(n_703), .S(n_702));
   FA_X1 i_378 (.A(n_698), .B(n_681), .CI(n_700), .CO(n_705), .S(n_704));
   FA_X1 i_379 (.A(n_702), .B(n_683), .CI(n_704), .CO(n_707), .S(n_706));
   HA_X1 i_380 (.A(n_685), .B(n_706), .CO(n_709), .S(n_708));
   XNOR2_X1 i_381 (.A(subRes3[42]), .B(subRes4[42]), .ZN(n_710));
   XNOR2_X1 i_382 (.A(n_710), .B(subRes5[42]), .ZN(n_711));
   INV_X1 i_383 (.A(n_711), .ZN(n_712));
   NAND3_X1 i_384 (.A1(n_714), .A2(n_716), .A3(n_717), .ZN(n_713));
   NAND2_X1 i_385 (.A1(subRes4[42]), .A2(n_715), .ZN(n_714));
   INV_X1 i_386 (.A(subRes3[42]), .ZN(n_715));
   NAND2_X1 i_387 (.A1(subRes5[42]), .A2(n_715), .ZN(n_716));
   NAND2_X1 i_388 (.A1(subRes5[42]), .A2(subRes4[42]), .ZN(n_717));
   FA_X1 i_389 (.A(subRes6[42]), .B(subRes7[42]), .CI(subRes8[42]), .CO(n_719), 
      .S(n_718));
   FA_X1 i_390 (.A(subRes9[42]), .B(subRes10[42]), .CI(subRes11[42]), .CO(n_721), 
      .S(n_720));
   FA_X1 i_391 (.A(subRes12[42]), .B(subRes13[42]), .CI(n_695), .CO(n_723), 
      .S(n_722));
   FA_X1 i_392 (.A(n_693), .B(n_691), .CI(n_689), .CO(n_725), .S(n_724));
   FA_X1 i_393 (.A(n_697), .B(n_722), .CI(n_720), .CO(n_727), .S(n_726));
   FA_X1 i_394 (.A(n_718), .B(n_712), .CI(n_724), .CO(n_729), .S(n_728));
   FA_X1 i_395 (.A(n_701), .B(n_699), .CI(n_703), .CO(n_731), .S(n_730));
   FA_X1 i_396 (.A(n_728), .B(n_726), .CI(n_730), .CO(n_733), .S(n_732));
   FA_X1 i_397 (.A(n_705), .B(n_732), .CI(n_707), .CO(n_735), .S(n_734));
   XNOR2_X1 i_398 (.A(subRes4[43]), .B(subRes5[43]), .ZN(n_736));
   OR2_X1 i_399 (.A1(subRes4[43]), .A2(subRes5[43]), .ZN(n_737));
   FA_X1 i_400 (.A(subRes6[43]), .B(subRes7[43]), .CI(subRes8[43]), .CO(n_739), 
      .S(n_738));
   FA_X1 i_401 (.A(subRes9[43]), .B(subRes10[43]), .CI(subRes11[43]), .CO(n_741), 
      .S(n_740));
   FA_X1 i_402 (.A(subRes12[43]), .B(subRes13[43]), .CI(n_721), .CO(n_743), 
      .S(n_742));
   FA_X1 i_403 (.A(n_719), .B(n_713), .CI(n_725), .CO(n_745), .S(n_744));
   FA_X1 i_404 (.A(n_723), .B(n_742), .CI(n_740), .CO(n_747), .S(n_746));
   FA_X1 i_405 (.A(n_738), .B(n_736), .CI(n_744), .CO(n_749), .S(n_748));
   FA_X1 i_406 (.A(n_727), .B(n_729), .CI(n_748), .CO(n_751), .S(n_750));
   FA_X1 i_407 (.A(n_746), .B(n_731), .CI(n_750), .CO(n_753), .S(n_752));
   HA_X1 i_408 (.A(n_733), .B(n_752), .CO(n_755), .S(n_754));
   XNOR2_X1 i_409 (.A(subRes4[44]), .B(subRes5[44]), .ZN(n_756));
   XNOR2_X1 i_410 (.A(n_756), .B(subRes6[44]), .ZN(n_757));
   INV_X1 i_411 (.A(n_757), .ZN(n_758));
   NAND3_X1 i_412 (.A1(n_760), .A2(n_762), .A3(n_763), .ZN(n_759));
   NAND2_X1 i_413 (.A1(subRes5[44]), .A2(n_761), .ZN(n_760));
   INV_X1 i_414 (.A(subRes4[44]), .ZN(n_761));
   NAND2_X1 i_415 (.A1(subRes6[44]), .A2(n_761), .ZN(n_762));
   NAND2_X1 i_416 (.A1(subRes6[44]), .A2(subRes5[44]), .ZN(n_763));
   FA_X1 i_417 (.A(subRes7[44]), .B(subRes8[44]), .CI(subRes9[44]), .CO(n_765), 
      .S(n_764));
   FA_X1 i_418 (.A(subRes10[44]), .B(subRes11[44]), .CI(subRes12[44]), .CO(n_767), 
      .S(n_766));
   FA_X1 i_419 (.A(subRes13[44]), .B(n_741), .CI(n_739), .CO(n_769), .S(n_768));
   FA_X1 i_420 (.A(n_737), .B(n_743), .CI(n_766), .CO(n_771), .S(n_770));
   FA_X1 i_421 (.A(n_764), .B(n_758), .CI(n_745), .CO(n_773), .S(n_772));
   FA_X1 i_422 (.A(n_768), .B(n_747), .CI(n_770), .CO(n_775), .S(n_774));
   FA_X1 i_423 (.A(n_749), .B(n_772), .CI(n_774), .CO(n_777), .S(n_776));
   FA_X1 i_424 (.A(n_751), .B(n_776), .CI(n_753), .CO(n_779), .S(n_778));
   XNOR2_X1 i_425 (.A(subRes5[45]), .B(subRes6[45]), .ZN(n_780));
   OR2_X1 i_426 (.A1(subRes5[45]), .A2(subRes6[45]), .ZN(n_781));
   FA_X1 i_427 (.A(subRes7[45]), .B(subRes8[45]), .CI(subRes9[45]), .CO(n_783), 
      .S(n_782));
   FA_X1 i_428 (.A(subRes10[45]), .B(subRes11[45]), .CI(subRes12[45]), .CO(n_785), 
      .S(n_784));
   FA_X1 i_429 (.A(subRes13[45]), .B(n_767), .CI(n_765), .CO(n_787), .S(n_786));
   FA_X1 i_430 (.A(n_759), .B(n_769), .CI(n_784), .CO(n_789), .S(n_788));
   FA_X1 i_431 (.A(n_782), .B(n_780), .CI(n_786), .CO(n_791), .S(n_790));
   FA_X1 i_432 (.A(n_771), .B(n_773), .CI(n_788), .CO(n_793), .S(n_792));
   FA_X1 i_433 (.A(n_790), .B(n_775), .CI(n_792), .CO(n_795), .S(n_794));
   HA_X1 i_434 (.A(n_777), .B(n_794), .CO(n_797), .S(n_796));
   XNOR2_X1 i_435 (.A(subRes5[46]), .B(subRes6[46]), .ZN(n_798));
   XNOR2_X1 i_436 (.A(n_798), .B(subRes7[46]), .ZN(n_799));
   INV_X1 i_437 (.A(n_799), .ZN(n_800));
   NAND3_X1 i_438 (.A1(n_802), .A2(n_804), .A3(n_805), .ZN(n_801));
   NAND2_X1 i_439 (.A1(subRes6[46]), .A2(n_803), .ZN(n_802));
   INV_X1 i_440 (.A(subRes5[46]), .ZN(n_803));
   NAND2_X1 i_441 (.A1(subRes7[46]), .A2(n_803), .ZN(n_804));
   NAND2_X1 i_442 (.A1(subRes7[46]), .A2(subRes6[46]), .ZN(n_805));
   FA_X1 i_443 (.A(subRes8[46]), .B(subRes9[46]), .CI(subRes10[46]), .CO(n_807), 
      .S(n_806));
   FA_X1 i_444 (.A(subRes11[46]), .B(subRes12[46]), .CI(subRes13[46]), .CO(n_809), 
      .S(n_808));
   FA_X1 i_445 (.A(n_785), .B(n_783), .CI(n_781), .CO(n_811), .S(n_810));
   FA_X1 i_446 (.A(n_787), .B(n_808), .CI(n_806), .CO(n_813), .S(n_812));
   FA_X1 i_447 (.A(n_800), .B(n_810), .CI(n_789), .CO(n_815), .S(n_814));
   FA_X1 i_448 (.A(n_791), .B(n_812), .CI(n_793), .CO(n_817), .S(n_816));
   FA_X1 i_449 (.A(n_814), .B(n_795), .CI(n_816), .CO(n_819), .S(n_818));
   XNOR2_X1 i_450 (.A(subRes6[47]), .B(subRes7[47]), .ZN(n_820));
   OR2_X1 i_451 (.A1(subRes6[47]), .A2(subRes7[47]), .ZN(n_821));
   FA_X1 i_452 (.A(subRes8[47]), .B(subRes9[47]), .CI(subRes10[47]), .CO(n_823), 
      .S(n_822));
   FA_X1 i_453 (.A(subRes11[47]), .B(subRes12[47]), .CI(subRes13[47]), .CO(n_825), 
      .S(n_824));
   FA_X1 i_454 (.A(n_809), .B(n_807), .CI(n_801), .CO(n_827), .S(n_826));
   FA_X1 i_455 (.A(n_811), .B(n_824), .CI(n_822), .CO(n_829), .S(n_828));
   FA_X1 i_456 (.A(n_820), .B(n_826), .CI(n_813), .CO(n_831), .S(n_830));
   FA_X1 i_457 (.A(n_815), .B(n_828), .CI(n_830), .CO(n_833), .S(n_832));
   HA_X1 i_458 (.A(n_817), .B(n_832), .CO(n_835), .S(n_834));
   XNOR2_X1 i_459 (.A(subRes6[48]), .B(subRes7[48]), .ZN(n_836));
   XNOR2_X1 i_460 (.A(n_836), .B(subRes8[48]), .ZN(n_837));
   INV_X1 i_461 (.A(n_837), .ZN(n_838));
   NAND3_X1 i_462 (.A1(n_840), .A2(n_842), .A3(n_843), .ZN(n_839));
   NAND2_X1 i_463 (.A1(subRes7[48]), .A2(n_841), .ZN(n_840));
   INV_X1 i_464 (.A(subRes6[48]), .ZN(n_841));
   NAND2_X1 i_465 (.A1(subRes8[48]), .A2(n_841), .ZN(n_842));
   NAND2_X1 i_466 (.A1(subRes8[48]), .A2(subRes7[48]), .ZN(n_843));
   FA_X1 i_467 (.A(subRes9[48]), .B(subRes10[48]), .CI(subRes11[48]), .CO(n_845), 
      .S(n_844));
   FA_X1 i_468 (.A(subRes12[48]), .B(subRes13[48]), .CI(n_825), .CO(n_847), 
      .S(n_846));
   FA_X1 i_469 (.A(n_823), .B(n_821), .CI(n_827), .CO(n_849), .S(n_848));
   FA_X1 i_470 (.A(n_846), .B(n_844), .CI(n_838), .CO(n_851), .S(n_850));
   FA_X1 i_471 (.A(n_848), .B(n_829), .CI(n_831), .CO(n_853), .S(n_852));
   FA_X1 i_472 (.A(n_850), .B(n_852), .CI(n_833), .CO(n_855), .S(n_854));
   XNOR2_X1 i_473 (.A(subRes7[49]), .B(subRes8[49]), .ZN(n_856));
   OR2_X1 i_474 (.A1(subRes7[49]), .A2(subRes8[49]), .ZN(n_857));
   FA_X1 i_475 (.A(subRes9[49]), .B(subRes10[49]), .CI(subRes11[49]), .CO(n_859), 
      .S(n_858));
   FA_X1 i_476 (.A(subRes12[49]), .B(subRes13[49]), .CI(n_845), .CO(n_861), 
      .S(n_860));
   FA_X1 i_477 (.A(n_839), .B(n_847), .CI(n_860), .CO(n_863), .S(n_862));
   FA_X1 i_478 (.A(n_858), .B(n_856), .CI(n_849), .CO(n_865), .S(n_864));
   FA_X1 i_479 (.A(n_851), .B(n_862), .CI(n_864), .CO(n_867), .S(n_866));
   HA_X1 i_480 (.A(n_853), .B(n_866), .CO(n_869), .S(n_868));
   XNOR2_X1 i_481 (.A(subRes7[50]), .B(subRes8[50]), .ZN(n_870));
   XNOR2_X1 i_482 (.A(n_870), .B(subRes9[50]), .ZN(n_871));
   INV_X1 i_483 (.A(n_871), .ZN(n_872));
   NAND3_X1 i_484 (.A1(n_874), .A2(n_876), .A3(n_877), .ZN(n_873));
   NAND2_X1 i_485 (.A1(subRes8[50]), .A2(n_875), .ZN(n_874));
   INV_X1 i_486 (.A(subRes7[50]), .ZN(n_875));
   NAND2_X1 i_487 (.A1(subRes9[50]), .A2(n_875), .ZN(n_876));
   NAND2_X1 i_488 (.A1(subRes9[50]), .A2(subRes8[50]), .ZN(n_877));
   FA_X1 i_489 (.A(subRes10[50]), .B(subRes11[50]), .CI(subRes12[50]), .CO(n_879), 
      .S(n_878));
   FA_X1 i_490 (.A(subRes13[50]), .B(n_859), .CI(n_857), .CO(n_881), .S(n_880));
   FA_X1 i_491 (.A(n_861), .B(n_878), .CI(n_872), .CO(n_883), .S(n_882));
   FA_X1 i_492 (.A(n_880), .B(n_863), .CI(n_865), .CO(n_885), .S(n_884));
   FA_X1 i_493 (.A(n_882), .B(n_884), .CI(n_867), .CO(n_887), .S(n_886));
   XNOR2_X1 i_494 (.A(subRes8[51]), .B(subRes9[51]), .ZN(n_888));
   OR2_X1 i_495 (.A1(subRes8[51]), .A2(subRes9[51]), .ZN(n_889));
   FA_X1 i_496 (.A(subRes10[51]), .B(subRes11[51]), .CI(subRes12[51]), .CO(n_891), 
      .S(n_890));
   FA_X1 i_497 (.A(subRes13[51]), .B(n_879), .CI(n_873), .CO(n_893), .S(n_892));
   FA_X1 i_498 (.A(n_881), .B(n_890), .CI(n_888), .CO(n_895), .S(n_894));
   FA_X1 i_499 (.A(n_892), .B(n_883), .CI(n_885), .CO(n_897), .S(n_896));
   HA_X1 i_500 (.A(n_894), .B(n_896), .CO(n_899), .S(n_898));
   XNOR2_X1 i_501 (.A(subRes8[52]), .B(subRes9[52]), .ZN(n_900));
   XNOR2_X1 i_502 (.A(n_900), .B(subRes10[52]), .ZN(n_901));
   INV_X1 i_503 (.A(n_901), .ZN(n_902));
   NAND3_X1 i_504 (.A1(n_904), .A2(n_906), .A3(n_907), .ZN(n_903));
   NAND2_X1 i_505 (.A1(subRes9[52]), .A2(n_905), .ZN(n_904));
   INV_X1 i_506 (.A(subRes8[52]), .ZN(n_905));
   NAND2_X1 i_507 (.A1(subRes10[52]), .A2(n_905), .ZN(n_906));
   NAND2_X1 i_508 (.A1(subRes10[52]), .A2(subRes9[52]), .ZN(n_907));
   FA_X1 i_509 (.A(subRes11[52]), .B(subRes12[52]), .CI(subRes13[52]), .CO(n_909), 
      .S(n_908));
   FA_X1 i_510 (.A(n_891), .B(n_889), .CI(n_893), .CO(n_911), .S(n_910));
   FA_X1 i_511 (.A(n_908), .B(n_902), .CI(n_910), .CO(n_913), .S(n_912));
   FA_X1 i_512 (.A(n_895), .B(n_912), .CI(n_897), .CO(n_915), .S(n_914));
   XNOR2_X1 i_513 (.A(subRes9[53]), .B(subRes10[53]), .ZN(n_916));
   OR2_X1 i_514 (.A1(subRes9[53]), .A2(subRes10[53]), .ZN(n_917));
   FA_X1 i_515 (.A(subRes11[53]), .B(subRes12[53]), .CI(subRes13[53]), .CO(n_919), 
      .S(n_918));
   FA_X1 i_516 (.A(n_909), .B(n_903), .CI(n_918), .CO(n_921), .S(n_920));
   FA_X1 i_517 (.A(n_916), .B(n_911), .CI(n_920), .CO(n_923), .S(n_922));
   HA_X1 i_518 (.A(n_913), .B(n_922), .CO(n_925), .S(n_924));
   XNOR2_X1 i_519 (.A(subRes9[54]), .B(subRes10[54]), .ZN(n_926));
   XNOR2_X1 i_520 (.A(n_926), .B(subRes11[54]), .ZN(n_927));
   INV_X1 i_521 (.A(n_927), .ZN(n_928));
   NAND3_X1 i_522 (.A1(n_930), .A2(n_932), .A3(n_933), .ZN(n_929));
   NAND2_X1 i_523 (.A1(subRes10[54]), .A2(n_931), .ZN(n_930));
   INV_X1 i_524 (.A(subRes9[54]), .ZN(n_931));
   NAND2_X1 i_525 (.A1(subRes11[54]), .A2(n_931), .ZN(n_932));
   NAND2_X1 i_526 (.A1(subRes11[54]), .A2(subRes10[54]), .ZN(n_933));
   FA_X1 i_527 (.A(subRes12[54]), .B(subRes13[54]), .CI(n_919), .CO(n_935), 
      .S(n_934));
   FA_X1 i_528 (.A(n_917), .B(n_934), .CI(n_928), .CO(n_937), .S(n_936));
   FA_X1 i_529 (.A(n_921), .B(n_923), .CI(n_936), .CO(n_939), .S(n_938));
   XNOR2_X1 i_530 (.A(subRes10[55]), .B(subRes11[55]), .ZN(n_940));
   OR2_X1 i_531 (.A1(subRes10[55]), .A2(subRes11[55]), .ZN(n_941));
   FA_X1 i_532 (.A(subRes12[55]), .B(subRes13[55]), .CI(n_929), .CO(n_943), 
      .S(n_942));
   FA_X1 i_533 (.A(n_935), .B(n_942), .CI(n_940), .CO(n_945), .S(n_944));
   HA_X1 i_534 (.A(n_937), .B(n_944), .CO(n_947), .S(n_946));
   XNOR2_X1 i_535 (.A(subRes10[56]), .B(subRes11[56]), .ZN(n_948));
   XNOR2_X1 i_536 (.A(n_948), .B(subRes12[56]), .ZN(n_949));
   INV_X1 i_537 (.A(n_949), .ZN(n_950));
   NAND3_X1 i_538 (.A1(n_952), .A2(n_954), .A3(n_955), .ZN(n_951));
   NAND2_X1 i_539 (.A1(subRes11[56]), .A2(n_953), .ZN(n_952));
   INV_X1 i_540 (.A(subRes10[56]), .ZN(n_953));
   NAND2_X1 i_541 (.A1(subRes12[56]), .A2(n_953), .ZN(n_954));
   NAND2_X1 i_542 (.A1(subRes12[56]), .A2(subRes11[56]), .ZN(n_955));
   FA_X1 i_543 (.A(subRes13[56]), .B(n_941), .CI(n_943), .CO(n_957), .S(n_956));
   FA_X1 i_544 (.A(n_950), .B(n_956), .CI(n_945), .CO(n_959), .S(n_958));
   XNOR2_X1 i_545 (.A(subRes11[57]), .B(subRes12[57]), .ZN(n_960));
   OR2_X1 i_546 (.A1(subRes11[57]), .A2(subRes12[57]), .ZN(n_961));
   FA_X1 i_547 (.A(subRes13[57]), .B(n_951), .CI(n_960), .CO(n_963), .S(n_962));
   HA_X1 i_548 (.A(n_957), .B(n_962), .CO(n_965), .S(n_964));
   XNOR2_X1 i_549 (.A(subRes11[58]), .B(subRes12[58]), .ZN(n_966));
   XNOR2_X1 i_550 (.A(n_966), .B(subRes13[58]), .ZN(n_967));
   INV_X1 i_551 (.A(n_967), .ZN(n_968));
   NAND3_X1 i_552 (.A1(n_970), .A2(n_972), .A3(n_973), .ZN(n_969));
   NAND2_X1 i_553 (.A1(subRes12[58]), .A2(n_971), .ZN(n_970));
   INV_X1 i_554 (.A(subRes11[58]), .ZN(n_971));
   NAND2_X1 i_555 (.A1(subRes13[58]), .A2(n_971), .ZN(n_972));
   NAND2_X1 i_556 (.A1(subRes13[58]), .A2(subRes12[58]), .ZN(n_973));
   FA_X1 i_557 (.A(n_961), .B(n_968), .CI(n_963), .CO(n_975), .S(n_974));
   XNOR2_X1 i_558 (.A(subRes12[59]), .B(subRes13[59]), .ZN(n_976));
   OR2_X1 i_559 (.A1(subRes12[59]), .A2(subRes13[59]), .ZN(n_977));
   HA_X1 i_560 (.A(n_969), .B(n_976), .CO(n_979), .S(n_978));
   XNOR2_X1 i_561 (.A(subRes12[60]), .B(subRes13[60]), .ZN(n_980));
   XNOR2_X1 i_562 (.A(n_980), .B(n_977), .ZN(n_981));
   INV_X1 i_563 (.A(n_981), .ZN(n_982));
   NAND3_X1 i_564 (.A1(n_984), .A2(n_986), .A3(n_987), .ZN(n_983));
   NAND2_X1 i_565 (.A1(subRes13[60]), .A2(n_985), .ZN(n_984));
   INV_X1 i_566 (.A(subRes12[60]), .ZN(n_985));
   NAND2_X1 i_567 (.A1(n_977), .A2(n_985), .ZN(n_986));
   NAND2_X1 i_568 (.A1(n_977), .A2(subRes13[60]), .ZN(n_987));
   INV_X1 i_569 (.A(subRes13[61]), .ZN(n_988));
   HA_X1 i_570 (.A(subRes[2]), .B(subRes14[2]), .CO(n_989), .S(product_reg[2]));
   FA_X1 i_571 (.A(subRes[3]), .B(subRes14[3]), .CI(n_989), .CO(n_990), .S(
      product_reg[3]));
   FA_X1 i_572 (.A(subRes14[4]), .B(n_0), .CI(n_990), .CO(n_991), .S(
      product_reg[4]));
   FA_X1 i_573 (.A(n_1), .B(n_2), .CI(n_991), .CO(n_992), .S(product_reg[5]));
   FA_X1 i_574 (.A(n_6), .B(n_4), .CI(n_992), .CO(n_993), .S(product_reg[6]));
   FA_X1 i_575 (.A(n_8), .B(n_10), .CI(n_993), .CO(n_994), .S(product_reg[7]));
   FA_X1 i_576 (.A(n_12), .B(n_16), .CI(n_994), .CO(n_995), .S(product_reg[8]));
   FA_X1 i_577 (.A(n_17), .B(n_22), .CI(n_995), .CO(n_996), .S(product_reg[9]));
   FA_X1 i_578 (.A(n_28), .B(n_30), .CI(n_996), .CO(n_997), .S(product_reg[10]));
   FA_X1 i_579 (.A(n_31), .B(n_38), .CI(n_997), .CO(n_998), .S(product_reg[11]));
   FA_X1 i_580 (.A(n_46), .B(n_48), .CI(n_998), .CO(n_999), .S(product_reg[12]));
   FA_X1 i_581 (.A(n_49), .B(n_58), .CI(n_999), .CO(n_1000), .S(product_reg[13]));
   FA_X1 i_582 (.A(n_59), .B(n_70), .CI(n_1000), .CO(n_1001), .S(product_reg[14]));
   FA_X1 i_583 (.A(n_71), .B(n_82), .CI(n_1001), .CO(n_1002), .S(product_reg[15]));
   FA_X1 i_584 (.A(n_83), .B(n_96), .CI(n_1002), .CO(n_1003), .S(product_reg[16]));
   FA_X1 i_585 (.A(n_97), .B(n_110), .CI(n_1003), .CO(n_1004), .S(
      product_reg[17]));
   FA_X1 i_586 (.A(n_111), .B(n_126), .CI(n_1004), .CO(n_1005), .S(
      product_reg[18]));
   FA_X1 i_587 (.A(n_127), .B(n_142), .CI(n_1005), .CO(n_1006), .S(
      product_reg[19]));
   FA_X1 i_588 (.A(n_143), .B(n_160), .CI(n_1006), .CO(n_1007), .S(
      product_reg[20]));
   FA_X1 i_589 (.A(n_161), .B(n_178), .CI(n_1007), .CO(n_1008), .S(
      product_reg[21]));
   FA_X1 i_590 (.A(n_179), .B(n_198), .CI(n_1008), .CO(n_1009), .S(
      product_reg[22]));
   FA_X1 i_591 (.A(n_199), .B(n_218), .CI(n_1009), .CO(n_1010), .S(
      product_reg[23]));
   FA_X1 i_592 (.A(n_219), .B(n_240), .CI(n_1010), .CO(n_1011), .S(
      product_reg[24]));
   FA_X1 i_593 (.A(n_241), .B(n_262), .CI(n_1011), .CO(n_1012), .S(
      product_reg[25]));
   FA_X1 i_594 (.A(n_263), .B(n_286), .CI(n_1012), .CO(n_1013), .S(
      product_reg[26]));
   FA_X1 i_595 (.A(n_287), .B(n_310), .CI(n_1013), .CO(n_1014), .S(
      product_reg[27]));
   FA_X1 i_596 (.A(n_311), .B(n_336), .CI(n_1014), .CO(n_1015), .S(
      product_reg[28]));
   FA_X1 i_597 (.A(n_337), .B(n_362), .CI(n_1015), .CO(n_1016), .S(
      product_reg[29]));
   FA_X1 i_598 (.A(n_363), .B(n_390), .CI(n_1016), .CO(n_1017), .S(
      product_reg[30]));
   FA_X1 i_599 (.A(n_391), .B(n_418), .CI(n_1017), .CO(n_1018), .S(
      product_reg[31]));
   FA_X1 i_600 (.A(n_419), .B(n_454), .CI(n_1018), .CO(n_1019), .S(
      product_reg[32]));
   FA_X1 i_601 (.A(n_455), .B(n_484), .CI(n_1019), .CO(n_1020), .S(
      product_reg[33]));
   FA_X1 i_602 (.A(n_485), .B(n_518), .CI(n_1020), .CO(n_1021), .S(
      product_reg[34]));
   FA_X1 i_603 (.A(n_519), .B(n_546), .CI(n_1021), .CO(n_1022), .S(
      product_reg[35]));
   FA_X1 i_604 (.A(n_547), .B(n_578), .CI(n_1022), .CO(n_1023), .S(
      product_reg[36]));
   FA_X1 i_605 (.A(n_579), .B(n_604), .CI(n_1023), .CO(n_1024), .S(
      product_reg[37]));
   FA_X1 i_606 (.A(n_605), .B(n_634), .CI(n_1024), .CO(n_1025), .S(
      product_reg[38]));
   FA_X1 i_607 (.A(n_635), .B(n_658), .CI(n_1025), .CO(n_1026), .S(
      product_reg[39]));
   FA_X1 i_608 (.A(n_659), .B(n_686), .CI(n_1026), .CO(n_1027), .S(
      product_reg[40]));
   FA_X1 i_609 (.A(n_687), .B(n_708), .CI(n_1027), .CO(n_1028), .S(
      product_reg[41]));
   FA_X1 i_610 (.A(n_709), .B(n_734), .CI(n_1028), .CO(n_1029), .S(
      product_reg[42]));
   FA_X1 i_611 (.A(n_735), .B(n_754), .CI(n_1029), .CO(n_1030), .S(
      product_reg[43]));
   FA_X1 i_612 (.A(n_755), .B(n_778), .CI(n_1030), .CO(n_1031), .S(
      product_reg[44]));
   FA_X1 i_613 (.A(n_779), .B(n_796), .CI(n_1031), .CO(n_1032), .S(
      product_reg[45]));
   FA_X1 i_614 (.A(n_797), .B(n_818), .CI(n_1032), .CO(n_1033), .S(
      product_reg[46]));
   FA_X1 i_615 (.A(n_819), .B(n_834), .CI(n_1033), .CO(n_1034), .S(
      product_reg[47]));
   FA_X1 i_616 (.A(n_835), .B(n_854), .CI(n_1034), .CO(n_1035), .S(
      product_reg[48]));
   FA_X1 i_617 (.A(n_855), .B(n_868), .CI(n_1035), .CO(n_1036), .S(
      product_reg[49]));
   FA_X1 i_618 (.A(n_869), .B(n_886), .CI(n_1036), .CO(n_1037), .S(
      product_reg[50]));
   FA_X1 i_619 (.A(n_887), .B(n_898), .CI(n_1037), .CO(n_1038), .S(
      product_reg[51]));
   FA_X1 i_620 (.A(n_899), .B(n_914), .CI(n_1038), .CO(n_1039), .S(
      product_reg[52]));
   FA_X1 i_621 (.A(n_915), .B(n_924), .CI(n_1039), .CO(n_1040), .S(
      product_reg[53]));
   FA_X1 i_622 (.A(n_925), .B(n_938), .CI(n_1040), .CO(n_1041), .S(
      product_reg[54]));
   FA_X1 i_623 (.A(n_939), .B(n_946), .CI(n_1041), .CO(n_1042), .S(
      product_reg[55]));
   FA_X1 i_624 (.A(n_947), .B(n_958), .CI(n_1042), .CO(n_1043), .S(
      product_reg[56]));
   FA_X1 i_625 (.A(n_959), .B(n_964), .CI(n_1043), .CO(n_1044), .S(
      product_reg[57]));
   FA_X1 i_626 (.A(n_965), .B(n_974), .CI(n_1044), .CO(n_1045), .S(
      product_reg[58]));
   FA_X1 i_627 (.A(n_978), .B(n_975), .CI(n_1045), .CO(n_1046), .S(
      product_reg[59]));
   FA_X1 i_628 (.A(n_982), .B(n_979), .CI(n_1046), .CO(n_1047), .S(
      product_reg[60]));
   FA_X1 i_629 (.A(n_988), .B(n_983), .CI(n_1047), .CO(n_1048), .S(
      product_reg[61]));
   XNOR2_X1 i_630 (.A(subRes13[62]), .B(subRes13[61]), .ZN(n_1049));
   XNOR2_X1 i_631 (.A(n_1049), .B(n_1048), .ZN(n_1050));
   INV_X1 i_632 (.A(n_1050), .ZN(product_reg[62]));
   NAND3_X1 i_633 (.A1(n_1052), .A2(n_1054), .A3(n_1055), .ZN(n_1051));
   NAND2_X1 i_634 (.A1(subRes13[61]), .A2(n_1053), .ZN(n_1052));
   INV_X1 i_635 (.A(subRes13[62]), .ZN(n_1053));
   NAND2_X1 i_636 (.A1(n_1048), .A2(n_1053), .ZN(n_1054));
   NAND2_X1 i_637 (.A1(n_1048), .A2(subRes13[61]), .ZN(n_1055));
   INV_X1 i_638 (.A(n_1051), .ZN(product_reg[63]));
endmodule

module Radix4BoothMultiplier(multiplicand, multiplier, product);
   input [31:0]multiplicand;
   input [31:0]multiplier;
   output [63:0]product;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_2_0;
   wire n_2_1;
   wire n_2_2;
   wire n_2_3;
   wire n_2_4;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire n_2_8;
   wire n_3_0;
   wire n_3_1;
   wire n_3_2;
   wire n_3_3;
   wire n_3_4;
   wire n_3_5;
   wire n_3_6;
   wire n_3_7;
   wire n_3_8;
   wire n_4_0;
   wire n_4_1;
   wire n_4_2;
   wire n_4_3;
   wire n_4_4;
   wire n_4_5;
   wire n_4_6;
   wire n_4_7;
   wire n_4_8;
   wire n_5_0;
   wire n_5_1;
   wire n_5_2;
   wire n_5_3;
   wire n_5_4;
   wire n_5_5;
   wire n_5_6;
   wire n_5_7;
   wire n_5_8;
   wire n_6_0;
   wire n_6_1;
   wire n_6_2;
   wire n_6_3;
   wire n_6_4;
   wire n_6_5;
   wire n_6_6;
   wire n_6_7;
   wire n_6_8;
   wire n_7_0;
   wire n_7_1;
   wire n_7_2;
   wire n_7_3;
   wire n_7_4;
   wire n_7_5;
   wire n_7_6;
   wire n_7_7;
   wire n_7_8;
   wire n_8_0;
   wire n_8_1;
   wire n_8_2;
   wire n_8_3;
   wire n_8_4;
   wire n_8_5;
   wire n_8_6;
   wire n_8_7;
   wire n_8_8;
   wire n_9_0;
   wire n_9_1;
   wire n_9_2;
   wire n_9_3;
   wire n_9_4;
   wire n_9_5;
   wire n_9_6;
   wire n_9_7;
   wire n_9_8;
   wire n_10_0;
   wire n_10_1;
   wire n_10_2;
   wire n_10_3;
   wire n_10_4;
   wire n_10_5;
   wire n_10_6;
   wire n_10_7;
   wire n_10_8;
   wire n_11_0;
   wire n_11_1;
   wire n_11_2;
   wire n_11_3;
   wire n_11_4;
   wire n_11_5;
   wire n_11_6;
   wire n_11_7;
   wire n_11_8;
   wire n_12_0;
   wire n_12_1;
   wire n_12_2;
   wire n_12_3;
   wire n_12_4;
   wire n_12_5;
   wire n_12_6;
   wire n_12_7;
   wire n_12_8;
   wire n_13_0;
   wire n_13_1;
   wire n_13_2;
   wire n_13_3;
   wire n_13_4;
   wire n_13_5;
   wire n_13_6;
   wire n_13_7;
   wire n_13_8;
   wire n_14_0;
   wire n_14_1;
   wire n_14_2;
   wire n_14_3;
   wire n_14_4;
   wire n_14_5;
   wire n_14_6;
   wire n_14_7;
   wire n_14_8;
   wire n_15_0;
   wire n_15_1;
   wire n_15_2;
   wire n_17_0;
   wire n_17_1;
   wire n_18_0;
   wire n_18_1;
   wire n_18_2;
   wire n_18_3;
   wire n_18_4;
   wire n_18_5;
   wire n_18_6;
   wire n_18_7;
   wire n_18_8;
   wire n_18_9;
   wire n_18_10;
   wire n_18_11;
   wire n_18_12;
   wire n_18_13;
   wire n_18_14;
   wire n_18_15;
   wire n_18_16;
   wire n_18_17;
   wire n_18_18;
   wire n_18_19;
   wire n_18_20;
   wire n_18_21;
   wire n_18_22;
   wire n_18_23;
   wire n_18_24;
   wire n_18_25;
   wire n_18_26;
   wire n_18_27;
   wire n_18_28;
   wire n_18_29;
   wire n_18_30;
   wire n_18_31;
   wire n_18_32;
   wire n_18_33;
   wire n_18_34;
   wire n_18_35;
   wire n_18_36;
   wire n_18_37;
   wire n_18_38;
   wire n_18_39;
   wire n_18_40;
   wire n_18_41;
   wire n_18_42;
   wire n_18_43;
   wire n_18_44;
   wire n_18_45;
   wire n_18_46;
   wire n_18_47;
   wire n_18_48;
   wire n_18_49;
   wire n_18_50;
   wire n_18_51;
   wire n_18_52;
   wire n_18_53;
   wire n_18_54;
   wire n_18_55;
   wire n_18_56;
   wire n_18_57;
   wire n_18_58;
   wire n_18_59;
   wire n_18_60;
   wire n_18_61;
   wire n_18_62;
   wire n_18_63;
   wire n_18_64;
   wire n_18_65;
   wire n_18_66;
   wire n_18_67;
   wire n_18_68;
   wire n_18_69;
   wire n_18_70;
   wire n_18_71;
   wire n_18_72;
   wire n_18_73;
   wire n_18_74;
   wire n_18_75;
   wire n_18_76;
   wire n_18_77;
   wire n_18_78;
   wire n_18_79;
   wire n_18_80;
   wire n_18_81;
   wire n_18_82;
   wire n_18_83;
   wire n_18_84;
   wire n_18_85;
   wire n_18_86;
   wire n_18_87;
   wire n_18_88;
   wire n_18_89;
   wire n_18_90;
   wire n_18_91;
   wire n_18_92;
   wire n_18_93;
   wire n_18_94;
   wire n_18_95;
   wire n_18_96;
   wire n_18_97;
   wire n_18_98;
   wire n_18_99;
   wire n_18_100;
   wire n_18_101;
   wire n_18_102;
   wire n_18_103;
   wire n_18_104;
   wire n_18_105;
   wire n_18_106;
   wire n_18_107;
   wire n_18_108;
   wire n_18_109;
   wire n_18_110;
   wire n_18_111;
   wire n_18_112;
   wire n_18_113;
   wire n_18_114;
   wire n_18_115;
   wire n_18_116;
   wire n_18_117;
   wire n_18_118;
   wire n_18_119;
   wire n_18_120;
   wire n_18_121;
   wire n_18_122;
   wire n_18_123;
   wire n_18_124;
   wire n_18_125;
   wire n_18_126;
   wire n_19_0;
   wire n_19_1;
   wire n_20_0;
   wire n_20_1;
   wire n_20_2;
   wire n_20_3;
   wire n_20_4;
   wire n_20_5;
   wire n_20_6;
   wire n_20_7;
   wire n_20_8;
   wire n_20_9;
   wire n_20_10;
   wire n_20_11;
   wire n_20_12;
   wire n_20_13;
   wire n_20_14;
   wire n_20_15;
   wire n_20_16;
   wire n_20_17;
   wire n_20_18;
   wire n_20_19;
   wire n_20_20;
   wire n_20_21;
   wire n_20_22;
   wire n_20_23;
   wire n_20_24;
   wire n_20_25;
   wire n_20_26;
   wire n_20_27;
   wire n_20_28;
   wire n_20_29;
   wire n_20_30;
   wire n_20_31;
   wire n_20_32;
   wire n_20_33;
   wire n_20_34;
   wire n_20_35;
   wire n_20_36;
   wire n_20_37;
   wire n_20_38;
   wire n_20_39;
   wire n_20_40;
   wire n_20_41;
   wire n_20_42;
   wire n_20_43;
   wire n_20_44;
   wire n_20_45;
   wire n_20_46;
   wire n_20_47;
   wire n_20_48;
   wire n_20_49;
   wire n_20_50;
   wire n_20_51;
   wire n_20_52;
   wire n_20_53;
   wire n_20_54;
   wire n_20_55;
   wire n_20_56;
   wire n_20_57;
   wire n_20_58;
   wire n_20_59;
   wire n_20_60;
   wire n_20_61;
   wire n_20_62;
   wire n_20_63;
   wire n_20_64;
   wire n_20_65;
   wire n_20_66;
   wire n_20_67;
   wire n_20_68;
   wire n_20_69;
   wire n_20_70;
   wire n_20_71;
   wire n_20_72;
   wire n_20_73;
   wire n_20_74;
   wire n_20_75;
   wire n_20_76;
   wire n_20_77;
   wire n_20_78;
   wire n_20_79;
   wire n_20_80;
   wire n_20_81;
   wire n_20_82;
   wire n_20_83;
   wire n_20_84;
   wire n_20_85;
   wire n_20_86;
   wire n_20_87;
   wire n_20_88;
   wire n_20_89;
   wire n_20_90;
   wire n_20_91;
   wire n_20_92;
   wire n_20_93;
   wire n_20_94;
   wire n_20_95;
   wire n_20_96;
   wire n_20_97;
   wire n_20_98;
   wire n_20_99;
   wire n_20_100;
   wire n_20_101;
   wire n_20_102;
   wire n_20_103;
   wire n_20_104;
   wire n_20_105;
   wire n_20_106;
   wire n_20_107;
   wire n_20_108;
   wire n_20_109;
   wire n_20_110;
   wire n_20_111;
   wire n_20_112;
   wire n_20_113;
   wire n_20_114;
   wire n_20_115;
   wire n_20_116;
   wire n_20_117;
   wire n_20_118;
   wire n_20_119;
   wire n_20_120;
   wire n_20_121;
   wire n_20_122;
   wire n_20_123;
   wire n_20_124;
   wire n_20_125;
   wire n_20_126;
   wire n_21_0;
   wire n_21_1;
   wire n_22_0;
   wire n_22_1;
   wire n_22_2;
   wire n_22_3;
   wire n_22_4;
   wire n_22_5;
   wire n_22_6;
   wire n_22_7;
   wire n_22_8;
   wire n_22_9;
   wire n_22_10;
   wire n_22_11;
   wire n_22_12;
   wire n_22_13;
   wire n_22_14;
   wire n_22_15;
   wire n_22_16;
   wire n_22_17;
   wire n_22_18;
   wire n_22_19;
   wire n_22_20;
   wire n_22_21;
   wire n_22_22;
   wire n_22_23;
   wire n_22_24;
   wire n_22_25;
   wire n_22_26;
   wire n_22_27;
   wire n_22_28;
   wire n_22_29;
   wire n_22_30;
   wire n_22_31;
   wire n_22_32;
   wire n_22_33;
   wire n_22_34;
   wire n_22_35;
   wire n_22_36;
   wire n_22_37;
   wire n_22_38;
   wire n_22_39;
   wire n_22_40;
   wire n_22_41;
   wire n_22_42;
   wire n_22_43;
   wire n_22_44;
   wire n_22_45;
   wire n_22_46;
   wire n_22_47;
   wire n_22_48;
   wire n_22_49;
   wire n_22_50;
   wire n_22_51;
   wire n_22_52;
   wire n_22_53;
   wire n_22_54;
   wire n_22_55;
   wire n_22_56;
   wire n_22_57;
   wire n_22_58;
   wire n_22_59;
   wire n_22_60;
   wire n_22_61;
   wire n_22_62;
   wire n_22_63;
   wire n_22_64;
   wire n_22_65;
   wire n_22_66;
   wire n_22_67;
   wire n_22_68;
   wire n_22_69;
   wire n_22_70;
   wire n_22_71;
   wire n_22_72;
   wire n_22_73;
   wire n_22_74;
   wire n_22_75;
   wire n_22_76;
   wire n_22_77;
   wire n_22_78;
   wire n_22_79;
   wire n_22_80;
   wire n_22_81;
   wire n_22_82;
   wire n_22_83;
   wire n_22_84;
   wire n_22_85;
   wire n_22_86;
   wire n_22_87;
   wire n_22_88;
   wire n_22_89;
   wire n_22_90;
   wire n_22_91;
   wire n_22_92;
   wire n_22_93;
   wire n_22_94;
   wire n_22_95;
   wire n_22_96;
   wire n_22_97;
   wire n_22_98;
   wire n_22_99;
   wire n_22_100;
   wire n_22_101;
   wire n_22_102;
   wire n_22_103;
   wire n_22_104;
   wire n_22_105;
   wire n_22_106;
   wire n_22_107;
   wire n_22_108;
   wire n_22_109;
   wire n_22_110;
   wire n_22_111;
   wire n_22_112;
   wire n_22_113;
   wire n_22_114;
   wire n_22_115;
   wire n_22_116;
   wire n_22_117;
   wire n_22_118;
   wire n_22_119;
   wire n_22_120;
   wire n_22_121;
   wire n_22_122;
   wire n_22_123;
   wire n_22_124;
   wire n_22_125;
   wire n_22_126;
   wire n_23_0;
   wire n_23_1;
   wire n_24_0;
   wire n_24_1;
   wire n_24_2;
   wire n_24_3;
   wire n_24_4;
   wire n_24_5;
   wire n_24_6;
   wire n_24_7;
   wire n_24_8;
   wire n_24_9;
   wire n_24_10;
   wire n_24_11;
   wire n_24_12;
   wire n_24_13;
   wire n_24_14;
   wire n_24_15;
   wire n_24_16;
   wire n_24_17;
   wire n_24_18;
   wire n_24_19;
   wire n_24_20;
   wire n_24_21;
   wire n_24_22;
   wire n_24_23;
   wire n_24_24;
   wire n_24_25;
   wire n_24_26;
   wire n_24_27;
   wire n_24_28;
   wire n_24_29;
   wire n_24_30;
   wire n_24_31;
   wire n_24_32;
   wire n_24_33;
   wire n_24_34;
   wire n_24_35;
   wire n_24_36;
   wire n_24_37;
   wire n_24_38;
   wire n_24_39;
   wire n_24_40;
   wire n_24_41;
   wire n_24_42;
   wire n_24_43;
   wire n_24_44;
   wire n_24_45;
   wire n_24_46;
   wire n_24_47;
   wire n_24_48;
   wire n_24_49;
   wire n_24_50;
   wire n_24_51;
   wire n_24_52;
   wire n_24_53;
   wire n_24_54;
   wire n_24_55;
   wire n_24_56;
   wire n_24_57;
   wire n_24_58;
   wire n_24_59;
   wire n_24_60;
   wire n_24_61;
   wire n_24_62;
   wire n_24_63;
   wire n_24_64;
   wire n_24_65;
   wire n_24_66;
   wire n_24_67;
   wire n_24_68;
   wire n_24_69;
   wire n_24_70;
   wire n_24_71;
   wire n_24_72;
   wire n_24_73;
   wire n_24_74;
   wire n_24_75;
   wire n_24_76;
   wire n_24_77;
   wire n_24_78;
   wire n_24_79;
   wire n_24_80;
   wire n_24_81;
   wire n_24_82;
   wire n_24_83;
   wire n_24_84;
   wire n_24_85;
   wire n_24_86;
   wire n_24_87;
   wire n_24_88;
   wire n_24_89;
   wire n_24_90;
   wire n_24_91;
   wire n_24_92;
   wire n_24_93;
   wire n_24_94;
   wire n_24_95;
   wire n_24_96;
   wire n_24_97;
   wire n_24_98;
   wire n_24_99;
   wire n_24_100;
   wire n_24_101;
   wire n_24_102;
   wire n_24_103;
   wire n_24_104;
   wire n_24_105;
   wire n_24_106;
   wire n_24_107;
   wire n_24_108;
   wire n_24_109;
   wire n_24_110;
   wire n_24_111;
   wire n_24_112;
   wire n_24_113;
   wire n_24_114;
   wire n_24_115;
   wire n_24_116;
   wire n_24_117;
   wire n_24_118;
   wire n_24_119;
   wire n_24_120;
   wire n_24_121;
   wire n_24_122;
   wire n_24_123;
   wire n_24_124;
   wire n_24_125;
   wire n_24_126;
   wire n_25_0;
   wire n_25_1;
   wire n_26_0;
   wire n_26_1;
   wire n_26_2;
   wire n_26_3;
   wire n_26_4;
   wire n_26_5;
   wire n_26_6;
   wire n_26_7;
   wire n_26_8;
   wire n_26_9;
   wire n_26_10;
   wire n_26_11;
   wire n_26_12;
   wire n_26_13;
   wire n_26_14;
   wire n_26_15;
   wire n_26_16;
   wire n_26_17;
   wire n_26_18;
   wire n_26_19;
   wire n_26_20;
   wire n_26_21;
   wire n_26_22;
   wire n_26_23;
   wire n_26_24;
   wire n_26_25;
   wire n_26_26;
   wire n_26_27;
   wire n_26_28;
   wire n_26_29;
   wire n_26_30;
   wire n_26_31;
   wire n_26_32;
   wire n_26_33;
   wire n_26_34;
   wire n_26_35;
   wire n_26_36;
   wire n_26_37;
   wire n_26_38;
   wire n_26_39;
   wire n_26_40;
   wire n_26_41;
   wire n_26_42;
   wire n_26_43;
   wire n_26_44;
   wire n_26_45;
   wire n_26_46;
   wire n_26_47;
   wire n_26_48;
   wire n_26_49;
   wire n_26_50;
   wire n_26_51;
   wire n_26_52;
   wire n_26_53;
   wire n_26_54;
   wire n_26_55;
   wire n_26_56;
   wire n_26_57;
   wire n_26_58;
   wire n_26_59;
   wire n_26_60;
   wire n_26_61;
   wire n_26_62;
   wire n_26_63;
   wire n_26_64;
   wire n_26_65;
   wire n_26_66;
   wire n_26_67;
   wire n_26_68;
   wire n_26_69;
   wire n_26_70;
   wire n_26_71;
   wire n_26_72;
   wire n_26_73;
   wire n_26_74;
   wire n_26_75;
   wire n_26_76;
   wire n_26_77;
   wire n_26_78;
   wire n_26_79;
   wire n_26_80;
   wire n_26_81;
   wire n_26_82;
   wire n_26_83;
   wire n_26_84;
   wire n_26_85;
   wire n_26_86;
   wire n_26_87;
   wire n_26_88;
   wire n_26_89;
   wire n_26_90;
   wire n_26_91;
   wire n_26_92;
   wire n_26_93;
   wire n_26_94;
   wire n_26_95;
   wire n_26_96;
   wire n_26_97;
   wire n_26_98;
   wire n_26_99;
   wire n_26_100;
   wire n_26_101;
   wire n_26_102;
   wire n_26_103;
   wire n_26_104;
   wire n_26_105;
   wire n_26_106;
   wire n_26_107;
   wire n_26_108;
   wire n_26_109;
   wire n_26_110;
   wire n_26_111;
   wire n_26_112;
   wire n_26_113;
   wire n_26_114;
   wire n_26_115;
   wire n_26_116;
   wire n_26_117;
   wire n_26_118;
   wire n_26_119;
   wire n_26_120;
   wire n_26_121;
   wire n_26_122;
   wire n_26_123;
   wire n_26_124;
   wire n_26_125;
   wire n_26_126;
   wire n_27_0;
   wire n_27_1;
   wire n_28_0;
   wire n_28_1;
   wire n_28_2;
   wire n_28_3;
   wire n_28_4;
   wire n_28_5;
   wire n_28_6;
   wire n_28_7;
   wire n_28_8;
   wire n_28_9;
   wire n_28_10;
   wire n_28_11;
   wire n_28_12;
   wire n_28_13;
   wire n_28_14;
   wire n_28_15;
   wire n_28_16;
   wire n_28_17;
   wire n_28_18;
   wire n_28_19;
   wire n_28_20;
   wire n_28_21;
   wire n_28_22;
   wire n_28_23;
   wire n_28_24;
   wire n_28_25;
   wire n_28_26;
   wire n_28_27;
   wire n_28_28;
   wire n_28_29;
   wire n_28_30;
   wire n_28_31;
   wire n_28_32;
   wire n_28_33;
   wire n_28_34;
   wire n_28_35;
   wire n_28_36;
   wire n_28_37;
   wire n_28_38;
   wire n_28_39;
   wire n_28_40;
   wire n_28_41;
   wire n_28_42;
   wire n_28_43;
   wire n_28_44;
   wire n_28_45;
   wire n_28_46;
   wire n_28_47;
   wire n_28_48;
   wire n_28_49;
   wire n_28_50;
   wire n_28_51;
   wire n_28_52;
   wire n_28_53;
   wire n_28_54;
   wire n_28_55;
   wire n_28_56;
   wire n_28_57;
   wire n_28_58;
   wire n_28_59;
   wire n_28_60;
   wire n_28_61;
   wire n_28_62;
   wire n_28_63;
   wire n_28_64;
   wire n_28_65;
   wire n_28_66;
   wire n_28_67;
   wire n_28_68;
   wire n_28_69;
   wire n_28_70;
   wire n_28_71;
   wire n_28_72;
   wire n_28_73;
   wire n_28_74;
   wire n_28_75;
   wire n_28_76;
   wire n_28_77;
   wire n_28_78;
   wire n_28_79;
   wire n_28_80;
   wire n_28_81;
   wire n_28_82;
   wire n_28_83;
   wire n_28_84;
   wire n_28_85;
   wire n_28_86;
   wire n_28_87;
   wire n_28_88;
   wire n_28_89;
   wire n_28_90;
   wire n_28_91;
   wire n_28_92;
   wire n_28_93;
   wire n_28_94;
   wire n_28_95;
   wire n_28_96;
   wire n_28_97;
   wire n_28_98;
   wire n_28_99;
   wire n_28_100;
   wire n_28_101;
   wire n_28_102;
   wire n_28_103;
   wire n_28_104;
   wire n_28_105;
   wire n_28_106;
   wire n_28_107;
   wire n_28_108;
   wire n_28_109;
   wire n_28_110;
   wire n_28_111;
   wire n_28_112;
   wire n_28_113;
   wire n_28_114;
   wire n_28_115;
   wire n_28_116;
   wire n_28_117;
   wire n_28_118;
   wire n_28_119;
   wire n_28_120;
   wire n_28_121;
   wire n_28_122;
   wire n_28_123;
   wire n_28_124;
   wire n_28_125;
   wire n_28_126;
   wire n_29_0;
   wire n_29_1;
   wire n_30_0;
   wire n_30_1;
   wire n_30_2;
   wire n_30_3;
   wire n_30_4;
   wire n_30_5;
   wire n_30_6;
   wire n_30_7;
   wire n_30_8;
   wire n_30_9;
   wire n_30_10;
   wire n_30_11;
   wire n_30_12;
   wire n_30_13;
   wire n_30_14;
   wire n_30_15;
   wire n_30_16;
   wire n_30_17;
   wire n_30_18;
   wire n_30_19;
   wire n_30_20;
   wire n_30_21;
   wire n_30_22;
   wire n_30_23;
   wire n_30_24;
   wire n_30_25;
   wire n_30_26;
   wire n_30_27;
   wire n_30_28;
   wire n_30_29;
   wire n_30_30;
   wire n_30_31;
   wire n_30_32;
   wire n_30_33;
   wire n_30_34;
   wire n_30_35;
   wire n_30_36;
   wire n_30_37;
   wire n_30_38;
   wire n_30_39;
   wire n_30_40;
   wire n_30_41;
   wire n_30_42;
   wire n_30_43;
   wire n_30_44;
   wire n_30_45;
   wire n_30_46;
   wire n_30_47;
   wire n_30_48;
   wire n_30_49;
   wire n_30_50;
   wire n_30_51;
   wire n_30_52;
   wire n_30_53;
   wire n_30_54;
   wire n_30_55;
   wire n_30_56;
   wire n_30_57;
   wire n_30_58;
   wire n_30_59;
   wire n_30_60;
   wire n_30_61;
   wire n_30_62;
   wire n_30_63;
   wire n_30_64;
   wire n_30_65;
   wire n_30_66;
   wire n_30_67;
   wire n_30_68;
   wire n_30_69;
   wire n_30_70;
   wire n_30_71;
   wire n_30_72;
   wire n_30_73;
   wire n_30_74;
   wire n_30_75;
   wire n_30_76;
   wire n_30_77;
   wire n_30_78;
   wire n_30_79;
   wire n_30_80;
   wire n_30_81;
   wire n_30_82;
   wire n_30_83;
   wire n_30_84;
   wire n_30_85;
   wire n_30_86;
   wire n_30_87;
   wire n_30_88;
   wire n_30_89;
   wire n_30_90;
   wire n_30_91;
   wire n_30_92;
   wire n_30_93;
   wire n_30_94;
   wire n_30_95;
   wire n_30_96;
   wire n_30_97;
   wire n_30_98;
   wire n_30_99;
   wire n_30_100;
   wire n_30_101;
   wire n_30_102;
   wire n_30_103;
   wire n_30_104;
   wire n_30_105;
   wire n_30_106;
   wire n_30_107;
   wire n_30_108;
   wire n_30_109;
   wire n_30_110;
   wire n_30_111;
   wire n_30_112;
   wire n_30_113;
   wire n_30_114;
   wire n_30_115;
   wire n_30_116;
   wire n_30_117;
   wire n_30_118;
   wire n_30_119;
   wire n_30_120;
   wire n_30_121;
   wire n_30_122;
   wire n_30_123;
   wire n_30_124;
   wire n_30_125;
   wire n_30_126;
   wire n_31_0;
   wire n_31_1;
   wire n_32_0;
   wire n_32_1;
   wire n_32_2;
   wire n_32_3;
   wire n_32_4;
   wire n_32_5;
   wire n_32_6;
   wire n_32_7;
   wire n_32_8;
   wire n_32_9;
   wire n_32_10;
   wire n_32_11;
   wire n_32_12;
   wire n_32_13;
   wire n_32_14;
   wire n_32_15;
   wire n_32_16;
   wire n_32_17;
   wire n_32_18;
   wire n_32_19;
   wire n_32_20;
   wire n_32_21;
   wire n_32_22;
   wire n_32_23;
   wire n_32_24;
   wire n_32_25;
   wire n_32_26;
   wire n_32_27;
   wire n_32_28;
   wire n_32_29;
   wire n_32_30;
   wire n_32_31;
   wire n_32_32;
   wire n_32_33;
   wire n_32_34;
   wire n_32_35;
   wire n_32_36;
   wire n_32_37;
   wire n_32_38;
   wire n_32_39;
   wire n_32_40;
   wire n_32_41;
   wire n_32_42;
   wire n_32_43;
   wire n_32_44;
   wire n_32_45;
   wire n_32_46;
   wire n_32_47;
   wire n_32_48;
   wire n_32_49;
   wire n_32_50;
   wire n_32_51;
   wire n_32_52;
   wire n_32_53;
   wire n_32_54;
   wire n_32_55;
   wire n_32_56;
   wire n_32_57;
   wire n_32_58;
   wire n_32_59;
   wire n_32_60;
   wire n_32_61;
   wire n_32_62;
   wire n_32_63;
   wire n_32_64;
   wire n_32_65;
   wire n_32_66;
   wire n_32_67;
   wire n_32_68;
   wire n_32_69;
   wire n_32_70;
   wire n_32_71;
   wire n_32_72;
   wire n_32_73;
   wire n_32_74;
   wire n_32_75;
   wire n_32_76;
   wire n_32_77;
   wire n_32_78;
   wire n_32_79;
   wire n_32_80;
   wire n_32_81;
   wire n_32_82;
   wire n_32_83;
   wire n_32_84;
   wire n_32_85;
   wire n_32_86;
   wire n_32_87;
   wire n_32_88;
   wire n_32_89;
   wire n_32_90;
   wire n_32_91;
   wire n_32_92;
   wire n_32_93;
   wire n_32_94;
   wire n_32_95;
   wire n_32_96;
   wire n_32_97;
   wire n_32_98;
   wire n_32_99;
   wire n_32_100;
   wire n_32_101;
   wire n_32_102;
   wire n_32_103;
   wire n_32_104;
   wire n_32_105;
   wire n_32_106;
   wire n_32_107;
   wire n_32_108;
   wire n_32_109;
   wire n_32_110;
   wire n_32_111;
   wire n_32_112;
   wire n_32_113;
   wire n_32_114;
   wire n_32_115;
   wire n_32_116;
   wire n_32_117;
   wire n_32_118;
   wire n_32_119;
   wire n_32_120;
   wire n_32_121;
   wire n_32_122;
   wire n_32_123;
   wire n_32_124;
   wire n_32_125;
   wire n_32_126;
   wire n_33_0;
   wire n_33_1;
   wire n_34_0;
   wire n_34_1;
   wire n_34_2;
   wire n_34_3;
   wire n_34_4;
   wire n_34_5;
   wire n_34_6;
   wire n_34_7;
   wire n_34_8;
   wire n_34_9;
   wire n_34_10;
   wire n_34_11;
   wire n_34_12;
   wire n_34_13;
   wire n_34_14;
   wire n_34_15;
   wire n_34_16;
   wire n_34_17;
   wire n_34_18;
   wire n_34_19;
   wire n_34_20;
   wire n_34_21;
   wire n_34_22;
   wire n_34_23;
   wire n_34_24;
   wire n_34_25;
   wire n_34_26;
   wire n_34_27;
   wire n_34_28;
   wire n_34_29;
   wire n_34_30;
   wire n_34_31;
   wire n_34_32;
   wire n_34_33;
   wire n_34_34;
   wire n_34_35;
   wire n_34_36;
   wire n_34_37;
   wire n_34_38;
   wire n_34_39;
   wire n_34_40;
   wire n_34_41;
   wire n_34_42;
   wire n_34_43;
   wire n_34_44;
   wire n_34_45;
   wire n_34_46;
   wire n_34_47;
   wire n_34_48;
   wire n_34_49;
   wire n_34_50;
   wire n_34_51;
   wire n_34_52;
   wire n_34_53;
   wire n_34_54;
   wire n_34_55;
   wire n_34_56;
   wire n_34_57;
   wire n_34_58;
   wire n_34_59;
   wire n_34_60;
   wire n_34_61;
   wire n_34_62;
   wire n_34_63;
   wire n_34_64;
   wire n_34_65;
   wire n_34_66;
   wire n_34_67;
   wire n_34_68;
   wire n_34_69;
   wire n_34_70;
   wire n_34_71;
   wire n_34_72;
   wire n_34_73;
   wire n_34_74;
   wire n_34_75;
   wire n_34_76;
   wire n_34_77;
   wire n_34_78;
   wire n_34_79;
   wire n_34_80;
   wire n_34_81;
   wire n_34_82;
   wire n_34_83;
   wire n_34_84;
   wire n_34_85;
   wire n_34_86;
   wire n_34_87;
   wire n_34_88;
   wire n_34_89;
   wire n_34_90;
   wire n_34_91;
   wire n_34_92;
   wire n_34_93;
   wire n_34_94;
   wire n_34_95;
   wire n_34_96;
   wire n_34_97;
   wire n_34_98;
   wire n_34_99;
   wire n_34_100;
   wire n_34_101;
   wire n_34_102;
   wire n_34_103;
   wire n_34_104;
   wire n_34_105;
   wire n_34_106;
   wire n_34_107;
   wire n_34_108;
   wire n_34_109;
   wire n_34_110;
   wire n_34_111;
   wire n_34_112;
   wire n_34_113;
   wire n_34_114;
   wire n_34_115;
   wire n_34_116;
   wire n_34_117;
   wire n_34_118;
   wire n_34_119;
   wire n_34_120;
   wire n_34_121;
   wire n_34_122;
   wire n_34_123;
   wire n_34_124;
   wire n_34_125;
   wire n_34_126;
   wire n_35_0;
   wire n_35_1;
   wire n_36_0;
   wire n_36_1;
   wire n_36_2;
   wire n_36_3;
   wire n_36_4;
   wire n_36_5;
   wire n_36_6;
   wire n_36_7;
   wire n_36_8;
   wire n_36_9;
   wire n_36_10;
   wire n_36_11;
   wire n_36_12;
   wire n_36_13;
   wire n_36_14;
   wire n_36_15;
   wire n_36_16;
   wire n_36_17;
   wire n_36_18;
   wire n_36_19;
   wire n_36_20;
   wire n_36_21;
   wire n_36_22;
   wire n_36_23;
   wire n_36_24;
   wire n_36_25;
   wire n_36_26;
   wire n_36_27;
   wire n_36_28;
   wire n_36_29;
   wire n_36_30;
   wire n_36_31;
   wire n_36_32;
   wire n_36_33;
   wire n_36_34;
   wire n_36_35;
   wire n_36_36;
   wire n_36_37;
   wire n_36_38;
   wire n_36_39;
   wire n_36_40;
   wire n_36_41;
   wire n_36_42;
   wire n_36_43;
   wire n_36_44;
   wire n_36_45;
   wire n_36_46;
   wire n_36_47;
   wire n_36_48;
   wire n_36_49;
   wire n_36_50;
   wire n_36_51;
   wire n_36_52;
   wire n_36_53;
   wire n_36_54;
   wire n_36_55;
   wire n_36_56;
   wire n_36_57;
   wire n_36_58;
   wire n_36_59;
   wire n_36_60;
   wire n_36_61;
   wire n_36_62;
   wire n_36_63;
   wire n_36_64;
   wire n_36_65;
   wire n_36_66;
   wire n_36_67;
   wire n_36_68;
   wire n_36_69;
   wire n_36_70;
   wire n_36_71;
   wire n_36_72;
   wire n_36_73;
   wire n_36_74;
   wire n_36_75;
   wire n_36_76;
   wire n_36_77;
   wire n_36_78;
   wire n_36_79;
   wire n_36_80;
   wire n_36_81;
   wire n_36_82;
   wire n_36_83;
   wire n_36_84;
   wire n_36_85;
   wire n_36_86;
   wire n_36_87;
   wire n_36_88;
   wire n_36_89;
   wire n_36_90;
   wire n_36_91;
   wire n_36_92;
   wire n_36_93;
   wire n_36_94;
   wire n_36_95;
   wire n_36_96;
   wire n_36_97;
   wire n_36_98;
   wire n_36_99;
   wire n_36_100;
   wire n_36_101;
   wire n_36_102;
   wire n_36_103;
   wire n_36_104;
   wire n_36_105;
   wire n_36_106;
   wire n_36_107;
   wire n_36_108;
   wire n_36_109;
   wire n_36_110;
   wire n_36_111;
   wire n_36_112;
   wire n_36_113;
   wire n_36_114;
   wire n_36_115;
   wire n_36_116;
   wire n_36_117;
   wire n_36_118;
   wire n_36_119;
   wire n_36_120;
   wire n_36_121;
   wire n_36_122;
   wire n_36_123;
   wire n_36_124;
   wire n_36_125;
   wire n_36_126;
   wire n_37_0;
   wire n_37_1;
   wire n_38_0;
   wire n_38_1;
   wire n_38_2;
   wire n_38_3;
   wire n_38_4;
   wire n_38_5;
   wire n_38_6;
   wire n_38_7;
   wire n_38_8;
   wire n_38_9;
   wire n_38_10;
   wire n_38_11;
   wire n_38_12;
   wire n_38_13;
   wire n_38_14;
   wire n_38_15;
   wire n_38_16;
   wire n_38_17;
   wire n_38_18;
   wire n_38_19;
   wire n_38_20;
   wire n_38_21;
   wire n_38_22;
   wire n_38_23;
   wire n_38_24;
   wire n_38_25;
   wire n_38_26;
   wire n_38_27;
   wire n_38_28;
   wire n_38_29;
   wire n_38_30;
   wire n_38_31;
   wire n_38_32;
   wire n_38_33;
   wire n_38_34;
   wire n_38_35;
   wire n_38_36;
   wire n_38_37;
   wire n_38_38;
   wire n_38_39;
   wire n_38_40;
   wire n_38_41;
   wire n_38_42;
   wire n_38_43;
   wire n_38_44;
   wire n_38_45;
   wire n_38_46;
   wire n_38_47;
   wire n_38_48;
   wire n_38_49;
   wire n_38_50;
   wire n_38_51;
   wire n_38_52;
   wire n_38_53;
   wire n_38_54;
   wire n_38_55;
   wire n_38_56;
   wire n_38_57;
   wire n_38_58;
   wire n_38_59;
   wire n_38_60;
   wire n_38_61;
   wire n_38_62;
   wire n_38_63;
   wire n_38_64;
   wire n_38_65;
   wire n_38_66;
   wire n_38_67;
   wire n_38_68;
   wire n_38_69;
   wire n_38_70;
   wire n_38_71;
   wire n_38_72;
   wire n_38_73;
   wire n_38_74;
   wire n_38_75;
   wire n_38_76;
   wire n_38_77;
   wire n_38_78;
   wire n_38_79;
   wire n_38_80;
   wire n_38_81;
   wire n_38_82;
   wire n_38_83;
   wire n_38_84;
   wire n_38_85;
   wire n_38_86;
   wire n_38_87;
   wire n_38_88;
   wire n_38_89;
   wire n_38_90;
   wire n_38_91;
   wire n_38_92;
   wire n_38_93;
   wire n_38_94;
   wire n_38_95;
   wire n_38_96;
   wire n_38_97;
   wire n_38_98;
   wire n_38_99;
   wire n_38_100;
   wire n_38_101;
   wire n_38_102;
   wire n_38_103;
   wire n_38_104;
   wire n_38_105;
   wire n_38_106;
   wire n_38_107;
   wire n_38_108;
   wire n_38_109;
   wire n_38_110;
   wire n_38_111;
   wire n_38_112;
   wire n_38_113;
   wire n_38_114;
   wire n_38_115;
   wire n_38_116;
   wire n_38_117;
   wire n_38_118;
   wire n_38_119;
   wire n_38_120;
   wire n_38_121;
   wire n_38_122;
   wire n_38_123;
   wire n_38_124;
   wire n_38_125;
   wire n_38_126;
   wire n_39_0;
   wire n_39_1;
   wire n_40_0;
   wire n_40_1;
   wire n_40_2;
   wire n_40_3;
   wire n_40_4;
   wire n_40_5;
   wire n_40_6;
   wire n_40_7;
   wire n_40_8;
   wire n_40_9;
   wire n_40_10;
   wire n_40_11;
   wire n_40_12;
   wire n_40_13;
   wire n_40_14;
   wire n_40_15;
   wire n_40_16;
   wire n_40_17;
   wire n_40_18;
   wire n_40_19;
   wire n_40_20;
   wire n_40_21;
   wire n_40_22;
   wire n_40_23;
   wire n_40_24;
   wire n_40_25;
   wire n_40_26;
   wire n_40_27;
   wire n_40_28;
   wire n_40_29;
   wire n_40_30;
   wire n_40_31;
   wire n_40_32;
   wire n_40_33;
   wire n_40_34;
   wire n_40_35;
   wire n_40_36;
   wire n_40_37;
   wire n_40_38;
   wire n_40_39;
   wire n_40_40;
   wire n_40_41;
   wire n_40_42;
   wire n_40_43;
   wire n_40_44;
   wire n_40_45;
   wire n_40_46;
   wire n_40_47;
   wire n_40_48;
   wire n_40_49;
   wire n_40_50;
   wire n_40_51;
   wire n_40_52;
   wire n_40_53;
   wire n_40_54;
   wire n_40_55;
   wire n_40_56;
   wire n_40_57;
   wire n_40_58;
   wire n_40_59;
   wire n_40_60;
   wire n_40_61;
   wire n_40_62;
   wire n_40_63;
   wire n_40_64;
   wire n_40_65;
   wire n_40_66;
   wire n_40_67;
   wire n_40_68;
   wire n_40_69;
   wire n_40_70;
   wire n_40_71;
   wire n_40_72;
   wire n_40_73;
   wire n_40_74;
   wire n_40_75;
   wire n_40_76;
   wire n_40_77;
   wire n_40_78;
   wire n_40_79;
   wire n_40_80;
   wire n_40_81;
   wire n_40_82;
   wire n_40_83;
   wire n_40_84;
   wire n_40_85;
   wire n_40_86;
   wire n_40_87;
   wire n_40_88;
   wire n_40_89;
   wire n_40_90;
   wire n_40_91;
   wire n_40_92;
   wire n_40_93;
   wire n_40_94;
   wire n_40_95;
   wire n_40_96;
   wire n_40_97;
   wire n_40_98;
   wire n_40_99;
   wire n_40_100;
   wire n_40_101;
   wire n_40_102;
   wire n_40_103;
   wire n_40_104;
   wire n_40_105;
   wire n_40_106;
   wire n_40_107;
   wire n_40_108;
   wire n_40_109;
   wire n_40_110;
   wire n_40_111;
   wire n_40_112;
   wire n_40_113;
   wire n_40_114;
   wire n_40_115;
   wire n_40_116;
   wire n_40_117;
   wire n_40_118;
   wire n_40_119;
   wire n_40_120;
   wire n_40_121;
   wire n_40_122;
   wire n_40_123;
   wire n_40_124;
   wire n_40_125;
   wire n_40_126;
   wire n_41_0;
   wire n_41_1;
   wire n_42_0;
   wire n_42_1;
   wire n_42_2;
   wire n_42_3;
   wire n_42_4;
   wire n_42_5;
   wire n_42_6;
   wire n_42_7;
   wire n_42_8;
   wire n_42_9;
   wire n_42_10;
   wire n_42_11;
   wire n_42_12;
   wire n_42_13;
   wire n_42_14;
   wire n_42_15;
   wire n_42_16;
   wire n_42_17;
   wire n_42_18;
   wire n_42_19;
   wire n_42_20;
   wire n_42_21;
   wire n_42_22;
   wire n_42_23;
   wire n_42_24;
   wire n_42_25;
   wire n_42_26;
   wire n_42_27;
   wire n_42_28;
   wire n_42_29;
   wire n_42_30;
   wire n_42_31;
   wire n_42_32;
   wire n_42_33;
   wire n_42_34;
   wire n_42_35;
   wire n_42_36;
   wire n_42_37;
   wire n_42_38;
   wire n_42_39;
   wire n_42_40;
   wire n_42_41;
   wire n_42_42;
   wire n_42_43;
   wire n_42_44;
   wire n_42_45;
   wire n_42_46;
   wire n_42_47;
   wire n_42_48;
   wire n_42_49;
   wire n_42_50;
   wire n_42_51;
   wire n_42_52;
   wire n_42_53;
   wire n_42_54;
   wire n_42_55;
   wire n_42_56;
   wire n_42_57;
   wire n_42_58;
   wire n_42_59;
   wire n_42_60;
   wire n_42_61;
   wire n_42_62;
   wire n_42_63;
   wire n_42_64;
   wire n_42_65;
   wire n_42_66;
   wire n_42_67;
   wire n_42_68;
   wire n_42_69;
   wire n_42_70;
   wire n_42_71;
   wire n_42_72;
   wire n_42_73;
   wire n_42_74;
   wire n_42_75;
   wire n_42_76;
   wire n_42_77;
   wire n_42_78;
   wire n_42_79;
   wire n_42_80;
   wire n_42_81;
   wire n_42_82;
   wire n_42_83;
   wire n_42_84;
   wire n_42_85;
   wire n_42_86;
   wire n_42_87;
   wire n_42_88;
   wire n_42_89;
   wire n_42_90;
   wire n_42_91;
   wire n_42_92;
   wire n_42_93;
   wire n_42_94;
   wire n_42_95;
   wire n_42_96;
   wire n_42_97;
   wire n_42_98;
   wire n_42_99;
   wire n_42_100;
   wire n_42_101;
   wire n_42_102;
   wire n_42_103;
   wire n_42_104;
   wire n_42_105;
   wire n_42_106;
   wire n_42_107;
   wire n_42_108;
   wire n_42_109;
   wire n_42_110;
   wire n_42_111;
   wire n_42_112;
   wire n_42_113;
   wire n_42_114;
   wire n_42_115;
   wire n_42_116;
   wire n_42_117;
   wire n_42_118;
   wire n_42_119;
   wire n_42_120;
   wire n_42_121;
   wire n_42_122;
   wire n_42_123;
   wire n_42_124;
   wire n_42_125;
   wire n_42_126;
   wire n_43_0;
   wire n_43_1;
   wire n_44_0;
   wire n_44_1;
   wire n_44_2;
   wire n_44_3;
   wire n_44_4;
   wire n_44_5;
   wire n_44_6;
   wire n_44_7;
   wire n_44_8;
   wire n_44_9;
   wire n_44_10;
   wire n_44_11;
   wire n_44_12;
   wire n_44_13;
   wire n_44_14;
   wire n_44_15;
   wire n_44_16;
   wire n_44_17;
   wire n_44_18;
   wire n_44_19;
   wire n_44_20;
   wire n_44_21;
   wire n_44_22;
   wire n_44_23;
   wire n_44_24;
   wire n_44_25;
   wire n_44_26;
   wire n_44_27;
   wire n_44_28;
   wire n_44_29;
   wire n_44_30;
   wire n_44_31;
   wire n_44_32;
   wire n_44_33;
   wire n_44_34;
   wire n_44_35;
   wire n_44_36;
   wire n_44_37;
   wire n_44_38;
   wire n_44_39;
   wire n_44_40;
   wire n_44_41;
   wire n_44_42;
   wire n_44_43;
   wire n_44_44;
   wire n_44_45;
   wire n_44_46;
   wire n_44_47;
   wire n_44_48;
   wire n_44_49;
   wire n_44_50;
   wire n_44_51;
   wire n_44_52;
   wire n_44_53;
   wire n_44_54;
   wire n_44_55;
   wire n_44_56;
   wire n_44_57;
   wire n_44_58;
   wire n_44_59;
   wire n_44_60;
   wire n_44_61;
   wire n_44_62;
   wire n_44_63;
   wire n_44_64;
   wire n_44_65;
   wire n_44_66;
   wire n_44_67;
   wire n_44_68;
   wire n_44_69;
   wire n_44_70;
   wire n_44_71;
   wire n_44_72;
   wire n_44_73;
   wire n_44_74;
   wire n_44_75;
   wire n_44_76;
   wire n_44_77;
   wire n_44_78;
   wire n_44_79;
   wire n_44_80;
   wire n_44_81;
   wire n_44_82;
   wire n_44_83;
   wire n_44_84;
   wire n_44_85;
   wire n_44_86;
   wire n_44_87;
   wire n_44_88;
   wire n_44_89;
   wire n_44_90;
   wire n_44_91;
   wire n_44_92;
   wire n_44_93;
   wire n_44_94;
   wire n_44_95;
   wire n_44_96;
   wire n_44_97;
   wire n_44_98;
   wire n_44_99;
   wire n_44_100;
   wire n_44_101;
   wire n_44_102;
   wire n_44_103;
   wire n_44_104;
   wire n_44_105;
   wire n_44_106;
   wire n_44_107;
   wire n_44_108;
   wire n_44_109;
   wire n_44_110;
   wire n_44_111;
   wire n_44_112;
   wire n_44_113;
   wire n_44_114;
   wire n_44_115;
   wire n_44_116;
   wire n_44_117;
   wire n_44_118;
   wire n_44_119;
   wire n_44_120;
   wire n_44_121;
   wire n_44_122;
   wire n_44_123;
   wire n_44_124;
   wire n_44_125;
   wire n_44_126;
   wire n_45_0;
   wire n_45_1;
   wire n_46_0;
   wire n_46_1;
   wire n_46_2;
   wire n_46_3;
   wire n_46_4;
   wire n_46_5;
   wire n_46_6;
   wire n_46_7;
   wire n_46_8;
   wire n_46_9;
   wire n_46_10;
   wire n_46_11;
   wire n_46_12;
   wire n_46_13;
   wire n_46_14;
   wire n_46_15;
   wire n_46_16;
   wire n_46_17;
   wire n_46_18;
   wire n_46_19;
   wire n_46_20;
   wire n_46_21;
   wire n_46_22;
   wire n_46_23;
   wire n_46_24;
   wire n_46_25;
   wire n_46_26;
   wire n_46_27;
   wire n_46_28;
   wire n_46_29;
   wire n_46_30;
   wire n_46_31;
   wire n_46_32;
   wire n_46_33;
   wire n_46_34;
   wire n_46_35;
   wire n_46_36;
   wire n_46_37;
   wire n_46_38;
   wire n_46_39;
   wire n_46_40;
   wire n_46_41;
   wire n_46_42;
   wire n_46_43;
   wire n_46_44;
   wire n_46_45;
   wire n_46_46;
   wire n_46_47;
   wire n_46_48;
   wire n_46_49;
   wire n_46_50;
   wire n_46_51;
   wire n_46_52;
   wire n_46_53;
   wire n_46_54;
   wire n_46_55;
   wire n_46_56;
   wire n_46_57;
   wire n_46_58;
   wire n_46_59;
   wire n_46_60;
   wire n_46_61;
   wire n_46_62;
   wire n_46_63;
   wire n_46_64;
   wire n_46_65;
   wire n_46_66;
   wire n_46_67;
   wire n_46_68;
   wire n_46_69;
   wire n_46_70;
   wire n_46_71;
   wire n_46_72;
   wire n_46_73;
   wire n_46_74;
   wire n_46_75;
   wire n_46_76;
   wire n_46_77;
   wire n_46_78;
   wire n_46_79;
   wire n_46_80;
   wire n_46_81;
   wire n_46_82;
   wire n_46_83;
   wire n_46_84;
   wire n_46_85;
   wire n_46_86;
   wire n_46_87;
   wire n_46_88;
   wire n_46_89;
   wire n_46_90;
   wire n_46_91;
   wire n_46_92;
   wire n_46_93;
   wire n_46_94;
   wire n_46_95;
   wire n_46_96;
   wire n_46_97;
   wire n_46_98;
   wire n_46_99;
   wire n_46_100;
   wire n_46_101;
   wire n_46_102;
   wire n_46_103;
   wire n_46_104;
   wire n_46_105;
   wire n_46_106;
   wire n_46_107;
   wire n_46_108;
   wire n_46_109;
   wire n_46_110;
   wire n_46_111;
   wire n_46_112;
   wire n_46_113;
   wire n_46_114;
   wire n_46_115;
   wire n_46_116;
   wire n_46_117;
   wire n_46_118;
   wire n_46_119;
   wire n_46_120;
   wire n_46_121;
   wire n_46_122;
   wire n_46_123;
   wire n_46_124;
   wire n_46_125;
   wire n_46_126;
   wire n_47_0;
   wire n_47_1;
   wire n_48_0;
   wire n_48_1;
   wire n_48_2;
   wire n_48_3;
   wire n_48_4;
   wire n_48_5;
   wire n_48_6;
   wire n_48_7;
   wire n_48_8;
   wire n_48_9;
   wire n_48_10;
   wire n_48_11;
   wire n_48_12;
   wire n_48_13;
   wire n_48_14;
   wire n_48_15;
   wire n_48_16;
   wire n_48_17;
   wire n_48_18;
   wire n_48_19;
   wire n_48_20;
   wire n_48_21;
   wire n_48_22;
   wire n_48_23;
   wire n_48_24;
   wire n_48_25;
   wire n_48_26;
   wire n_48_27;
   wire n_48_28;
   wire n_48_29;
   wire n_48_30;
   wire n_48_31;
   wire n_48_32;
   wire n_48_33;
   wire n_48_34;

   INV_X1 i_0_0 (.A(multiplier[2]), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(multiplier[1]), .ZN(n_0_1));
   OAI33_X1 i_0_2 (.A1(n_0_0), .A2(multiplier[1]), .A3(multiplier[3]), .B1(n_0_1), 
      .B2(multiplier[2]), .B3(multiplier[3]), .ZN(n_0_2));
   NAND3_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .A3(multiplier[3]), .ZN(n_0_3));
   OR3_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(multiplier[3]), .ZN(n_0_4));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0));
   INV_X1 i_0_6 (.A(n_0), .ZN(n_0_5));
   NAND3_X1 i_0_7 (.A1(n_0_1), .A2(multiplier[2]), .A3(multiplier[3]), .ZN(n_0_6));
   NAND3_X1 i_0_8 (.A1(n_0_0), .A2(multiplier[1]), .A3(multiplier[3]), .ZN(n_0_7));
   NAND4_X1 i_0_9 (.A1(n_0_2), .A2(n_0_5), .A3(n_0_6), .A4(n_0_7), .ZN(n_0_8));
   NAND3_X1 i_0_10 (.A1(n_0_8), .A2(n_0_6), .A3(n_0_7), .ZN(n_1));
   NAND3_X1 i_0_11 (.A1(n_0_3), .A2(n_0_6), .A3(n_0_7), .ZN(n_2));
   INV_X1 i_1_0 (.A(multiplier[4]), .ZN(n_1_0));
   INV_X1 i_1_1 (.A(multiplier[3]), .ZN(n_1_1));
   OAI33_X1 i_1_2 (.A1(n_1_0), .A2(multiplier[3]), .A3(multiplier[5]), .B1(n_1_1), 
      .B2(multiplier[4]), .B3(multiplier[5]), .ZN(n_1_2));
   NAND3_X1 i_1_3 (.A1(n_1_1), .A2(n_1_0), .A3(multiplier[5]), .ZN(n_1_3));
   OR3_X1 i_1_4 (.A1(n_1_0), .A2(n_1_1), .A3(multiplier[5]), .ZN(n_1_4));
   NAND2_X1 i_1_5 (.A1(n_1_3), .A2(n_1_4), .ZN(n_3));
   INV_X1 i_1_6 (.A(n_3), .ZN(n_1_5));
   NAND3_X1 i_1_7 (.A1(n_1_1), .A2(multiplier[4]), .A3(multiplier[5]), .ZN(n_1_6));
   NAND3_X1 i_1_8 (.A1(n_1_0), .A2(multiplier[3]), .A3(multiplier[5]), .ZN(n_1_7));
   NAND4_X1 i_1_9 (.A1(n_1_2), .A2(n_1_5), .A3(n_1_6), .A4(n_1_7), .ZN(n_1_8));
   NAND3_X1 i_1_10 (.A1(n_1_8), .A2(n_1_6), .A3(n_1_7), .ZN(n_4));
   NAND3_X1 i_1_11 (.A1(n_1_3), .A2(n_1_6), .A3(n_1_7), .ZN(n_5));
   INV_X1 i_2_0 (.A(multiplier[6]), .ZN(n_2_0));
   INV_X1 i_2_1 (.A(multiplier[5]), .ZN(n_2_1));
   OAI33_X1 i_2_2 (.A1(n_2_0), .A2(multiplier[5]), .A3(multiplier[7]), .B1(n_2_1), 
      .B2(multiplier[6]), .B3(multiplier[7]), .ZN(n_2_2));
   NAND3_X1 i_2_3 (.A1(n_2_1), .A2(n_2_0), .A3(multiplier[7]), .ZN(n_2_3));
   OR3_X1 i_2_4 (.A1(n_2_0), .A2(n_2_1), .A3(multiplier[7]), .ZN(n_2_4));
   NAND2_X1 i_2_5 (.A1(n_2_3), .A2(n_2_4), .ZN(n_6));
   INV_X1 i_2_6 (.A(n_6), .ZN(n_2_5));
   NAND3_X1 i_2_7 (.A1(n_2_1), .A2(multiplier[6]), .A3(multiplier[7]), .ZN(n_2_6));
   NAND3_X1 i_2_8 (.A1(n_2_0), .A2(multiplier[5]), .A3(multiplier[7]), .ZN(n_2_7));
   NAND4_X1 i_2_9 (.A1(n_2_2), .A2(n_2_5), .A3(n_2_6), .A4(n_2_7), .ZN(n_2_8));
   NAND3_X1 i_2_10 (.A1(n_2_8), .A2(n_2_6), .A3(n_2_7), .ZN(n_7));
   NAND3_X1 i_2_11 (.A1(n_2_3), .A2(n_2_6), .A3(n_2_7), .ZN(n_8));
   INV_X1 i_3_0 (.A(multiplier[8]), .ZN(n_3_0));
   INV_X1 i_3_1 (.A(multiplier[7]), .ZN(n_3_1));
   OAI33_X1 i_3_2 (.A1(n_3_0), .A2(multiplier[7]), .A3(multiplier[9]), .B1(n_3_1), 
      .B2(multiplier[8]), .B3(multiplier[9]), .ZN(n_3_2));
   NAND3_X1 i_3_3 (.A1(n_3_1), .A2(n_3_0), .A3(multiplier[9]), .ZN(n_3_3));
   OR3_X1 i_3_4 (.A1(n_3_0), .A2(n_3_1), .A3(multiplier[9]), .ZN(n_3_4));
   NAND2_X1 i_3_5 (.A1(n_3_3), .A2(n_3_4), .ZN(n_9));
   INV_X1 i_3_6 (.A(n_9), .ZN(n_3_5));
   NAND3_X1 i_3_7 (.A1(n_3_1), .A2(multiplier[8]), .A3(multiplier[9]), .ZN(n_3_6));
   NAND3_X1 i_3_8 (.A1(n_3_0), .A2(multiplier[7]), .A3(multiplier[9]), .ZN(n_3_7));
   NAND4_X1 i_3_9 (.A1(n_3_2), .A2(n_3_5), .A3(n_3_6), .A4(n_3_7), .ZN(n_3_8));
   NAND3_X1 i_3_10 (.A1(n_3_8), .A2(n_3_6), .A3(n_3_7), .ZN(n_10));
   NAND3_X1 i_3_11 (.A1(n_3_3), .A2(n_3_6), .A3(n_3_7), .ZN(n_11));
   INV_X1 i_4_0 (.A(multiplier[10]), .ZN(n_4_0));
   INV_X1 i_4_1 (.A(multiplier[9]), .ZN(n_4_1));
   OAI33_X1 i_4_2 (.A1(n_4_0), .A2(multiplier[9]), .A3(multiplier[11]), .B1(
      n_4_1), .B2(multiplier[10]), .B3(multiplier[11]), .ZN(n_4_2));
   NAND3_X1 i_4_3 (.A1(n_4_1), .A2(n_4_0), .A3(multiplier[11]), .ZN(n_4_3));
   OR3_X1 i_4_4 (.A1(n_4_0), .A2(n_4_1), .A3(multiplier[11]), .ZN(n_4_4));
   NAND2_X1 i_4_5 (.A1(n_4_3), .A2(n_4_4), .ZN(n_12));
   INV_X1 i_4_6 (.A(n_12), .ZN(n_4_5));
   NAND3_X1 i_4_7 (.A1(n_4_1), .A2(multiplier[10]), .A3(multiplier[11]), 
      .ZN(n_4_6));
   NAND3_X1 i_4_8 (.A1(n_4_0), .A2(multiplier[9]), .A3(multiplier[11]), .ZN(
      n_4_7));
   NAND4_X1 i_4_9 (.A1(n_4_2), .A2(n_4_5), .A3(n_4_6), .A4(n_4_7), .ZN(n_4_8));
   NAND3_X1 i_4_10 (.A1(n_4_8), .A2(n_4_6), .A3(n_4_7), .ZN(n_13));
   NAND3_X1 i_4_11 (.A1(n_4_3), .A2(n_4_6), .A3(n_4_7), .ZN(n_14));
   INV_X1 i_5_0 (.A(multiplier[12]), .ZN(n_5_0));
   INV_X1 i_5_1 (.A(multiplier[11]), .ZN(n_5_1));
   OAI33_X1 i_5_2 (.A1(n_5_0), .A2(multiplier[11]), .A3(multiplier[13]), 
      .B1(n_5_1), .B2(multiplier[12]), .B3(multiplier[13]), .ZN(n_5_2));
   NAND3_X1 i_5_3 (.A1(n_5_1), .A2(n_5_0), .A3(multiplier[13]), .ZN(n_5_3));
   OR3_X1 i_5_4 (.A1(n_5_0), .A2(n_5_1), .A3(multiplier[13]), .ZN(n_5_4));
   NAND2_X1 i_5_5 (.A1(n_5_3), .A2(n_5_4), .ZN(n_15));
   INV_X1 i_5_6 (.A(n_15), .ZN(n_5_5));
   NAND3_X1 i_5_7 (.A1(n_5_1), .A2(multiplier[12]), .A3(multiplier[13]), 
      .ZN(n_5_6));
   NAND3_X1 i_5_8 (.A1(n_5_0), .A2(multiplier[11]), .A3(multiplier[13]), 
      .ZN(n_5_7));
   NAND4_X1 i_5_9 (.A1(n_5_2), .A2(n_5_5), .A3(n_5_6), .A4(n_5_7), .ZN(n_5_8));
   NAND3_X1 i_5_10 (.A1(n_5_8), .A2(n_5_6), .A3(n_5_7), .ZN(n_16));
   NAND3_X1 i_5_11 (.A1(n_5_3), .A2(n_5_6), .A3(n_5_7), .ZN(n_17));
   INV_X1 i_6_0 (.A(multiplier[14]), .ZN(n_6_0));
   INV_X1 i_6_1 (.A(multiplier[13]), .ZN(n_6_1));
   OAI33_X1 i_6_2 (.A1(n_6_0), .A2(multiplier[13]), .A3(multiplier[15]), 
      .B1(n_6_1), .B2(multiplier[14]), .B3(multiplier[15]), .ZN(n_6_2));
   NAND3_X1 i_6_3 (.A1(n_6_1), .A2(n_6_0), .A3(multiplier[15]), .ZN(n_6_3));
   OR3_X1 i_6_4 (.A1(n_6_0), .A2(n_6_1), .A3(multiplier[15]), .ZN(n_6_4));
   NAND2_X1 i_6_5 (.A1(n_6_3), .A2(n_6_4), .ZN(n_18));
   INV_X1 i_6_6 (.A(n_18), .ZN(n_6_5));
   NAND3_X1 i_6_7 (.A1(n_6_1), .A2(multiplier[14]), .A3(multiplier[15]), 
      .ZN(n_6_6));
   NAND3_X1 i_6_8 (.A1(n_6_0), .A2(multiplier[13]), .A3(multiplier[15]), 
      .ZN(n_6_7));
   NAND4_X1 i_6_9 (.A1(n_6_2), .A2(n_6_5), .A3(n_6_6), .A4(n_6_7), .ZN(n_6_8));
   NAND3_X1 i_6_10 (.A1(n_6_8), .A2(n_6_6), .A3(n_6_7), .ZN(n_19));
   NAND3_X1 i_6_11 (.A1(n_6_3), .A2(n_6_6), .A3(n_6_7), .ZN(n_20));
   INV_X1 i_7_0 (.A(multiplier[16]), .ZN(n_7_0));
   INV_X1 i_7_1 (.A(multiplier[15]), .ZN(n_7_1));
   OAI33_X1 i_7_2 (.A1(n_7_0), .A2(multiplier[15]), .A3(multiplier[17]), 
      .B1(n_7_1), .B2(multiplier[16]), .B3(multiplier[17]), .ZN(n_7_2));
   NAND3_X1 i_7_3 (.A1(n_7_1), .A2(n_7_0), .A3(multiplier[17]), .ZN(n_7_3));
   OR3_X1 i_7_4 (.A1(n_7_0), .A2(n_7_1), .A3(multiplier[17]), .ZN(n_7_4));
   NAND2_X1 i_7_5 (.A1(n_7_3), .A2(n_7_4), .ZN(n_21));
   INV_X1 i_7_6 (.A(n_21), .ZN(n_7_5));
   NAND3_X1 i_7_7 (.A1(n_7_1), .A2(multiplier[16]), .A3(multiplier[17]), 
      .ZN(n_7_6));
   NAND3_X1 i_7_8 (.A1(n_7_0), .A2(multiplier[15]), .A3(multiplier[17]), 
      .ZN(n_7_7));
   NAND4_X1 i_7_9 (.A1(n_7_2), .A2(n_7_5), .A3(n_7_6), .A4(n_7_7), .ZN(n_7_8));
   NAND3_X1 i_7_10 (.A1(n_7_8), .A2(n_7_6), .A3(n_7_7), .ZN(n_22));
   NAND3_X1 i_7_11 (.A1(n_7_3), .A2(n_7_6), .A3(n_7_7), .ZN(n_23));
   INV_X1 i_8_0 (.A(multiplier[18]), .ZN(n_8_0));
   INV_X1 i_8_1 (.A(multiplier[17]), .ZN(n_8_1));
   OAI33_X1 i_8_2 (.A1(n_8_0), .A2(multiplier[17]), .A3(multiplier[19]), 
      .B1(n_8_1), .B2(multiplier[18]), .B3(multiplier[19]), .ZN(n_8_2));
   NAND3_X1 i_8_3 (.A1(n_8_1), .A2(n_8_0), .A3(multiplier[19]), .ZN(n_8_3));
   OR3_X1 i_8_4 (.A1(n_8_0), .A2(n_8_1), .A3(multiplier[19]), .ZN(n_8_4));
   NAND2_X1 i_8_5 (.A1(n_8_3), .A2(n_8_4), .ZN(n_24));
   INV_X1 i_8_6 (.A(n_24), .ZN(n_8_5));
   NAND3_X1 i_8_7 (.A1(n_8_1), .A2(multiplier[18]), .A3(multiplier[19]), 
      .ZN(n_8_6));
   NAND3_X1 i_8_8 (.A1(n_8_0), .A2(multiplier[17]), .A3(multiplier[19]), 
      .ZN(n_8_7));
   NAND4_X1 i_8_9 (.A1(n_8_2), .A2(n_8_5), .A3(n_8_6), .A4(n_8_7), .ZN(n_8_8));
   NAND3_X1 i_8_10 (.A1(n_8_8), .A2(n_8_6), .A3(n_8_7), .ZN(n_25));
   NAND3_X1 i_8_11 (.A1(n_8_3), .A2(n_8_6), .A3(n_8_7), .ZN(n_26));
   INV_X1 i_9_0 (.A(multiplier[20]), .ZN(n_9_0));
   INV_X1 i_9_1 (.A(multiplier[19]), .ZN(n_9_1));
   OAI33_X1 i_9_2 (.A1(n_9_0), .A2(multiplier[19]), .A3(multiplier[21]), 
      .B1(n_9_1), .B2(multiplier[20]), .B3(multiplier[21]), .ZN(n_9_2));
   NAND3_X1 i_9_3 (.A1(n_9_1), .A2(n_9_0), .A3(multiplier[21]), .ZN(n_9_3));
   OR3_X1 i_9_4 (.A1(n_9_0), .A2(n_9_1), .A3(multiplier[21]), .ZN(n_9_4));
   NAND2_X1 i_9_5 (.A1(n_9_3), .A2(n_9_4), .ZN(n_27));
   INV_X1 i_9_6 (.A(n_27), .ZN(n_9_5));
   NAND3_X1 i_9_7 (.A1(n_9_1), .A2(multiplier[20]), .A3(multiplier[21]), 
      .ZN(n_9_6));
   NAND3_X1 i_9_8 (.A1(n_9_0), .A2(multiplier[19]), .A3(multiplier[21]), 
      .ZN(n_9_7));
   NAND4_X1 i_9_9 (.A1(n_9_2), .A2(n_9_5), .A3(n_9_6), .A4(n_9_7), .ZN(n_9_8));
   NAND3_X1 i_9_10 (.A1(n_9_8), .A2(n_9_6), .A3(n_9_7), .ZN(n_28));
   NAND3_X1 i_9_11 (.A1(n_9_3), .A2(n_9_6), .A3(n_9_7), .ZN(n_29));
   INV_X1 i_10_0 (.A(multiplier[22]), .ZN(n_10_0));
   INV_X1 i_10_1 (.A(multiplier[21]), .ZN(n_10_1));
   OAI33_X1 i_10_2 (.A1(n_10_0), .A2(multiplier[21]), .A3(multiplier[23]), 
      .B1(n_10_1), .B2(multiplier[22]), .B3(multiplier[23]), .ZN(n_10_2));
   NAND3_X1 i_10_3 (.A1(n_10_1), .A2(n_10_0), .A3(multiplier[23]), .ZN(n_10_3));
   OR3_X1 i_10_4 (.A1(n_10_0), .A2(n_10_1), .A3(multiplier[23]), .ZN(n_10_4));
   NAND2_X1 i_10_5 (.A1(n_10_3), .A2(n_10_4), .ZN(n_30));
   INV_X1 i_10_6 (.A(n_30), .ZN(n_10_5));
   NAND3_X1 i_10_7 (.A1(n_10_1), .A2(multiplier[22]), .A3(multiplier[23]), 
      .ZN(n_10_6));
   NAND3_X1 i_10_8 (.A1(n_10_0), .A2(multiplier[21]), .A3(multiplier[23]), 
      .ZN(n_10_7));
   NAND4_X1 i_10_9 (.A1(n_10_2), .A2(n_10_5), .A3(n_10_6), .A4(n_10_7), .ZN(
      n_10_8));
   NAND3_X1 i_10_10 (.A1(n_10_8), .A2(n_10_6), .A3(n_10_7), .ZN(n_31));
   NAND3_X1 i_10_11 (.A1(n_10_3), .A2(n_10_6), .A3(n_10_7), .ZN(n_32));
   INV_X1 i_11_0 (.A(multiplier[24]), .ZN(n_11_0));
   INV_X1 i_11_1 (.A(multiplier[23]), .ZN(n_11_1));
   OAI33_X1 i_11_2 (.A1(n_11_0), .A2(multiplier[23]), .A3(multiplier[25]), 
      .B1(n_11_1), .B2(multiplier[24]), .B3(multiplier[25]), .ZN(n_11_2));
   NAND3_X1 i_11_3 (.A1(n_11_1), .A2(n_11_0), .A3(multiplier[25]), .ZN(n_11_3));
   OR3_X1 i_11_4 (.A1(n_11_0), .A2(n_11_1), .A3(multiplier[25]), .ZN(n_11_4));
   NAND2_X1 i_11_5 (.A1(n_11_3), .A2(n_11_4), .ZN(n_33));
   INV_X1 i_11_6 (.A(n_33), .ZN(n_11_5));
   NAND3_X1 i_11_7 (.A1(n_11_1), .A2(multiplier[24]), .A3(multiplier[25]), 
      .ZN(n_11_6));
   NAND3_X1 i_11_8 (.A1(n_11_0), .A2(multiplier[23]), .A3(multiplier[25]), 
      .ZN(n_11_7));
   NAND4_X1 i_11_9 (.A1(n_11_2), .A2(n_11_5), .A3(n_11_6), .A4(n_11_7), .ZN(
      n_11_8));
   NAND3_X1 i_11_10 (.A1(n_11_8), .A2(n_11_6), .A3(n_11_7), .ZN(n_34));
   NAND3_X1 i_11_11 (.A1(n_11_3), .A2(n_11_6), .A3(n_11_7), .ZN(n_35));
   INV_X1 i_12_0 (.A(multiplier[26]), .ZN(n_12_0));
   INV_X1 i_12_1 (.A(multiplier[25]), .ZN(n_12_1));
   OAI33_X1 i_12_2 (.A1(n_12_0), .A2(multiplier[25]), .A3(multiplier[27]), 
      .B1(n_12_1), .B2(multiplier[26]), .B3(multiplier[27]), .ZN(n_12_2));
   NAND3_X1 i_12_3 (.A1(n_12_1), .A2(n_12_0), .A3(multiplier[27]), .ZN(n_12_3));
   OR3_X1 i_12_4 (.A1(n_12_0), .A2(n_12_1), .A3(multiplier[27]), .ZN(n_12_4));
   NAND2_X1 i_12_5 (.A1(n_12_3), .A2(n_12_4), .ZN(n_36));
   INV_X1 i_12_6 (.A(n_36), .ZN(n_12_5));
   NAND3_X1 i_12_7 (.A1(n_12_1), .A2(multiplier[26]), .A3(multiplier[27]), 
      .ZN(n_12_6));
   NAND3_X1 i_12_8 (.A1(n_12_0), .A2(multiplier[25]), .A3(multiplier[27]), 
      .ZN(n_12_7));
   NAND4_X1 i_12_9 (.A1(n_12_2), .A2(n_12_5), .A3(n_12_6), .A4(n_12_7), .ZN(
      n_12_8));
   NAND3_X1 i_12_10 (.A1(n_12_8), .A2(n_12_6), .A3(n_12_7), .ZN(n_37));
   NAND3_X1 i_12_11 (.A1(n_12_3), .A2(n_12_6), .A3(n_12_7), .ZN(n_38));
   INV_X1 i_13_0 (.A(multiplier[28]), .ZN(n_13_0));
   INV_X1 i_13_1 (.A(multiplier[27]), .ZN(n_13_1));
   OAI33_X1 i_13_2 (.A1(n_13_0), .A2(multiplier[27]), .A3(multiplier[29]), 
      .B1(n_13_1), .B2(multiplier[28]), .B3(multiplier[29]), .ZN(n_13_2));
   NAND3_X1 i_13_3 (.A1(n_13_1), .A2(n_13_0), .A3(multiplier[29]), .ZN(n_13_3));
   OR3_X1 i_13_4 (.A1(n_13_0), .A2(n_13_1), .A3(multiplier[29]), .ZN(n_13_4));
   NAND2_X1 i_13_5 (.A1(n_13_3), .A2(n_13_4), .ZN(n_39));
   INV_X1 i_13_6 (.A(n_39), .ZN(n_13_5));
   NAND3_X1 i_13_7 (.A1(n_13_1), .A2(multiplier[28]), .A3(multiplier[29]), 
      .ZN(n_13_6));
   NAND3_X1 i_13_8 (.A1(n_13_0), .A2(multiplier[27]), .A3(multiplier[29]), 
      .ZN(n_13_7));
   NAND4_X1 i_13_9 (.A1(n_13_2), .A2(n_13_5), .A3(n_13_6), .A4(n_13_7), .ZN(
      n_13_8));
   NAND3_X1 i_13_10 (.A1(n_13_8), .A2(n_13_6), .A3(n_13_7), .ZN(n_40));
   NAND3_X1 i_13_11 (.A1(n_13_3), .A2(n_13_6), .A3(n_13_7), .ZN(n_41));
   INV_X1 i_14_0 (.A(multiplier[30]), .ZN(n_14_0));
   INV_X1 i_14_1 (.A(multiplier[29]), .ZN(n_14_1));
   OAI33_X1 i_14_2 (.A1(n_14_0), .A2(multiplier[29]), .A3(multiplier[31]), 
      .B1(n_14_1), .B2(multiplier[30]), .B3(multiplier[31]), .ZN(n_14_2));
   NAND3_X1 i_14_3 (.A1(n_14_1), .A2(n_14_0), .A3(multiplier[31]), .ZN(n_14_3));
   OR3_X1 i_14_4 (.A1(n_14_0), .A2(n_14_1), .A3(multiplier[31]), .ZN(n_14_4));
   NAND2_X1 i_14_5 (.A1(n_14_3), .A2(n_14_4), .ZN(n_42));
   INV_X1 i_14_6 (.A(n_42), .ZN(n_14_5));
   NAND3_X1 i_14_7 (.A1(n_14_1), .A2(multiplier[30]), .A3(multiplier[31]), 
      .ZN(n_14_6));
   NAND3_X1 i_14_8 (.A1(n_14_0), .A2(multiplier[29]), .A3(multiplier[31]), 
      .ZN(n_14_7));
   NAND4_X1 i_14_9 (.A1(n_14_2), .A2(n_14_5), .A3(n_14_6), .A4(n_14_7), .ZN(
      n_14_8));
   NAND3_X1 i_14_10 (.A1(n_14_8), .A2(n_14_6), .A3(n_14_7), .ZN(n_43));
   NAND3_X1 i_14_11 (.A1(n_14_3), .A2(n_14_6), .A3(n_14_7), .ZN(n_44));
   NAND2_X1 i_15_0 (.A1(multiplier[0]), .A2(multiplier[1]), .ZN(n_15_0));
   INV_X1 i_15_1 (.A(multiplier[0]), .ZN(n_15_1));
   OAI21_X1 i_15_2 (.A(n_15_0), .B1(n_15_1), .B2(multiplier[1]), .ZN(n_45));
   NAND2_X1 i_15_3 (.A1(n_15_1), .A2(multiplier[1]), .ZN(n_15_2));
   INV_X1 i_15_4 (.A(n_15_2), .ZN(n_46));
   NAND2_X1 i_15_5 (.A1(n_15_2), .A2(n_15_0), .ZN(n_47));
   datapath i_16 (.p_0({n_78, n_77, n_76, n_75, n_74, n_73, n_72, n_71, n_70, 
      n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, uc_0}), 
      .multiplicand(multiplicand));
   INV_X1 i_17_0 (.A(n_0), .ZN(n_17_0));
   AND3_X1 i_17_1 (.A1(n_17_0), .A2(n_1), .A3(n_2), .ZN(n_79));
   INV_X1 i_17_2 (.A(n_1), .ZN(n_17_1));
   AND3_X1 i_17_3 (.A1(n_17_1), .A2(n_0), .A3(n_2), .ZN(n_80));
   NOR3_X1 i_17_4 (.A1(n_17_1), .A2(n_0), .A3(n_2), .ZN(n_81));
   NOR3_X1 i_17_5 (.A1(n_17_0), .A2(n_1), .A3(n_2), .ZN(n_82));
   AOI22_X1 i_18_0 (.A1(n_81), .A2(multiplicand[0]), .B1(n_79), .B2(
      multiplicand[0]), .ZN(n_18_0));
   INV_X1 i_18_1 (.A(n_18_0), .ZN(n_83));
   NAND2_X1 i_18_2 (.A1(n_81), .A2(multiplicand[1]), .ZN(n_18_1));
   NAND2_X1 i_18_3 (.A1(n_79), .A2(n_48), .ZN(n_18_2));
   NAND2_X1 i_18_4 (.A1(n_80), .A2(multiplicand[0]), .ZN(n_18_3));
   NAND2_X1 i_18_5 (.A1(n_82), .A2(multiplicand[0]), .ZN(n_18_4));
   NAND4_X1 i_18_6 (.A1(n_18_1), .A2(n_18_2), .A3(n_18_3), .A4(n_18_4), .ZN(n_84));
   NAND2_X1 i_18_7 (.A1(n_81), .A2(multiplicand[2]), .ZN(n_18_5));
   NAND2_X1 i_18_8 (.A1(n_79), .A2(n_49), .ZN(n_18_6));
   NAND2_X1 i_18_9 (.A1(n_80), .A2(n_48), .ZN(n_18_7));
   NAND2_X1 i_18_10 (.A1(n_82), .A2(multiplicand[1]), .ZN(n_18_8));
   NAND4_X1 i_18_11 (.A1(n_18_5), .A2(n_18_6), .A3(n_18_7), .A4(n_18_8), 
      .ZN(n_85));
   NAND2_X1 i_18_12 (.A1(n_81), .A2(multiplicand[3]), .ZN(n_18_9));
   NAND2_X1 i_18_13 (.A1(n_79), .A2(n_50), .ZN(n_18_10));
   NAND2_X1 i_18_14 (.A1(n_80), .A2(n_49), .ZN(n_18_11));
   NAND2_X1 i_18_15 (.A1(n_82), .A2(multiplicand[2]), .ZN(n_18_12));
   NAND4_X1 i_18_16 (.A1(n_18_9), .A2(n_18_10), .A3(n_18_11), .A4(n_18_12), 
      .ZN(n_86));
   NAND2_X1 i_18_17 (.A1(n_81), .A2(multiplicand[4]), .ZN(n_18_13));
   NAND2_X1 i_18_18 (.A1(n_79), .A2(n_51), .ZN(n_18_14));
   NAND2_X1 i_18_19 (.A1(n_80), .A2(n_50), .ZN(n_18_15));
   NAND2_X1 i_18_20 (.A1(n_82), .A2(multiplicand[3]), .ZN(n_18_16));
   NAND4_X1 i_18_21 (.A1(n_18_13), .A2(n_18_14), .A3(n_18_15), .A4(n_18_16), 
      .ZN(n_87));
   NAND2_X1 i_18_22 (.A1(n_81), .A2(multiplicand[5]), .ZN(n_18_17));
   NAND2_X1 i_18_23 (.A1(n_79), .A2(n_52), .ZN(n_18_18));
   NAND2_X1 i_18_24 (.A1(n_80), .A2(n_51), .ZN(n_18_19));
   NAND2_X1 i_18_25 (.A1(n_82), .A2(multiplicand[4]), .ZN(n_18_20));
   NAND4_X1 i_18_26 (.A1(n_18_17), .A2(n_18_18), .A3(n_18_19), .A4(n_18_20), 
      .ZN(n_88));
   NAND2_X1 i_18_27 (.A1(n_81), .A2(multiplicand[6]), .ZN(n_18_21));
   NAND2_X1 i_18_28 (.A1(n_79), .A2(n_53), .ZN(n_18_22));
   NAND2_X1 i_18_29 (.A1(n_80), .A2(n_52), .ZN(n_18_23));
   NAND2_X1 i_18_30 (.A1(n_82), .A2(multiplicand[5]), .ZN(n_18_24));
   NAND4_X1 i_18_31 (.A1(n_18_21), .A2(n_18_22), .A3(n_18_23), .A4(n_18_24), 
      .ZN(n_89));
   NAND2_X1 i_18_32 (.A1(n_81), .A2(multiplicand[7]), .ZN(n_18_25));
   NAND2_X1 i_18_33 (.A1(n_79), .A2(n_54), .ZN(n_18_26));
   NAND2_X1 i_18_34 (.A1(n_80), .A2(n_53), .ZN(n_18_27));
   NAND2_X1 i_18_35 (.A1(n_82), .A2(multiplicand[6]), .ZN(n_18_28));
   NAND4_X1 i_18_36 (.A1(n_18_25), .A2(n_18_26), .A3(n_18_27), .A4(n_18_28), 
      .ZN(n_90));
   NAND2_X1 i_18_37 (.A1(n_81), .A2(multiplicand[8]), .ZN(n_18_29));
   NAND2_X1 i_18_38 (.A1(n_79), .A2(n_55), .ZN(n_18_30));
   NAND2_X1 i_18_39 (.A1(n_80), .A2(n_54), .ZN(n_18_31));
   NAND2_X1 i_18_40 (.A1(n_82), .A2(multiplicand[7]), .ZN(n_18_32));
   NAND4_X1 i_18_41 (.A1(n_18_29), .A2(n_18_30), .A3(n_18_31), .A4(n_18_32), 
      .ZN(n_91));
   NAND2_X1 i_18_42 (.A1(n_81), .A2(multiplicand[9]), .ZN(n_18_33));
   NAND2_X1 i_18_43 (.A1(n_79), .A2(n_56), .ZN(n_18_34));
   NAND2_X1 i_18_44 (.A1(n_80), .A2(n_55), .ZN(n_18_35));
   NAND2_X1 i_18_45 (.A1(n_82), .A2(multiplicand[8]), .ZN(n_18_36));
   NAND4_X1 i_18_46 (.A1(n_18_33), .A2(n_18_34), .A3(n_18_35), .A4(n_18_36), 
      .ZN(n_92));
   NAND2_X1 i_18_47 (.A1(n_81), .A2(multiplicand[10]), .ZN(n_18_37));
   NAND2_X1 i_18_48 (.A1(n_79), .A2(n_57), .ZN(n_18_38));
   NAND2_X1 i_18_49 (.A1(n_80), .A2(n_56), .ZN(n_18_39));
   NAND2_X1 i_18_50 (.A1(n_82), .A2(multiplicand[9]), .ZN(n_18_40));
   NAND4_X1 i_18_51 (.A1(n_18_37), .A2(n_18_38), .A3(n_18_39), .A4(n_18_40), 
      .ZN(n_93));
   NAND2_X1 i_18_52 (.A1(n_81), .A2(multiplicand[11]), .ZN(n_18_41));
   NAND2_X1 i_18_53 (.A1(n_79), .A2(n_58), .ZN(n_18_42));
   NAND2_X1 i_18_54 (.A1(n_80), .A2(n_57), .ZN(n_18_43));
   NAND2_X1 i_18_55 (.A1(n_82), .A2(multiplicand[10]), .ZN(n_18_44));
   NAND4_X1 i_18_56 (.A1(n_18_41), .A2(n_18_42), .A3(n_18_43), .A4(n_18_44), 
      .ZN(n_94));
   NAND2_X1 i_18_57 (.A1(n_81), .A2(multiplicand[12]), .ZN(n_18_45));
   NAND2_X1 i_18_58 (.A1(n_79), .A2(n_59), .ZN(n_18_46));
   NAND2_X1 i_18_59 (.A1(n_80), .A2(n_58), .ZN(n_18_47));
   NAND2_X1 i_18_60 (.A1(n_82), .A2(multiplicand[11]), .ZN(n_18_48));
   NAND4_X1 i_18_61 (.A1(n_18_45), .A2(n_18_46), .A3(n_18_47), .A4(n_18_48), 
      .ZN(n_95));
   NAND2_X1 i_18_62 (.A1(n_81), .A2(multiplicand[13]), .ZN(n_18_49));
   NAND2_X1 i_18_63 (.A1(n_79), .A2(n_60), .ZN(n_18_50));
   NAND2_X1 i_18_64 (.A1(n_80), .A2(n_59), .ZN(n_18_51));
   NAND2_X1 i_18_65 (.A1(n_82), .A2(multiplicand[12]), .ZN(n_18_52));
   NAND4_X1 i_18_66 (.A1(n_18_49), .A2(n_18_50), .A3(n_18_51), .A4(n_18_52), 
      .ZN(n_96));
   NAND2_X1 i_18_67 (.A1(n_81), .A2(multiplicand[14]), .ZN(n_18_53));
   NAND2_X1 i_18_68 (.A1(n_79), .A2(n_61), .ZN(n_18_54));
   NAND2_X1 i_18_69 (.A1(n_80), .A2(n_60), .ZN(n_18_55));
   NAND2_X1 i_18_70 (.A1(n_82), .A2(multiplicand[13]), .ZN(n_18_56));
   NAND4_X1 i_18_71 (.A1(n_18_53), .A2(n_18_54), .A3(n_18_55), .A4(n_18_56), 
      .ZN(n_97));
   NAND2_X1 i_18_72 (.A1(n_81), .A2(multiplicand[15]), .ZN(n_18_57));
   NAND2_X1 i_18_73 (.A1(n_79), .A2(n_62), .ZN(n_18_58));
   NAND2_X1 i_18_74 (.A1(n_80), .A2(n_61), .ZN(n_18_59));
   NAND2_X1 i_18_75 (.A1(n_82), .A2(multiplicand[14]), .ZN(n_18_60));
   NAND4_X1 i_18_76 (.A1(n_18_57), .A2(n_18_58), .A3(n_18_59), .A4(n_18_60), 
      .ZN(n_98));
   NAND2_X1 i_18_77 (.A1(n_81), .A2(multiplicand[16]), .ZN(n_18_61));
   NAND2_X1 i_18_78 (.A1(n_79), .A2(n_63), .ZN(n_18_62));
   NAND2_X1 i_18_79 (.A1(n_80), .A2(n_62), .ZN(n_18_63));
   NAND2_X1 i_18_80 (.A1(n_82), .A2(multiplicand[15]), .ZN(n_18_64));
   NAND4_X1 i_18_81 (.A1(n_18_61), .A2(n_18_62), .A3(n_18_63), .A4(n_18_64), 
      .ZN(n_99));
   NAND2_X1 i_18_82 (.A1(n_81), .A2(multiplicand[17]), .ZN(n_18_65));
   NAND2_X1 i_18_83 (.A1(n_79), .A2(n_64), .ZN(n_18_66));
   NAND2_X1 i_18_84 (.A1(n_80), .A2(n_63), .ZN(n_18_67));
   NAND2_X1 i_18_85 (.A1(n_82), .A2(multiplicand[16]), .ZN(n_18_68));
   NAND4_X1 i_18_86 (.A1(n_18_65), .A2(n_18_66), .A3(n_18_67), .A4(n_18_68), 
      .ZN(n_100));
   NAND2_X1 i_18_87 (.A1(n_81), .A2(multiplicand[18]), .ZN(n_18_69));
   NAND2_X1 i_18_88 (.A1(n_79), .A2(n_65), .ZN(n_18_70));
   NAND2_X1 i_18_89 (.A1(n_80), .A2(n_64), .ZN(n_18_71));
   NAND2_X1 i_18_90 (.A1(n_82), .A2(multiplicand[17]), .ZN(n_18_72));
   NAND4_X1 i_18_91 (.A1(n_18_69), .A2(n_18_70), .A3(n_18_71), .A4(n_18_72), 
      .ZN(n_101));
   NAND2_X1 i_18_92 (.A1(n_81), .A2(multiplicand[19]), .ZN(n_18_73));
   NAND2_X1 i_18_93 (.A1(n_79), .A2(n_66), .ZN(n_18_74));
   NAND2_X1 i_18_94 (.A1(n_80), .A2(n_65), .ZN(n_18_75));
   NAND2_X1 i_18_95 (.A1(n_82), .A2(multiplicand[18]), .ZN(n_18_76));
   NAND4_X1 i_18_96 (.A1(n_18_73), .A2(n_18_74), .A3(n_18_75), .A4(n_18_76), 
      .ZN(n_102));
   NAND2_X1 i_18_97 (.A1(n_81), .A2(multiplicand[20]), .ZN(n_18_77));
   NAND2_X1 i_18_98 (.A1(n_79), .A2(n_67), .ZN(n_18_78));
   NAND2_X1 i_18_99 (.A1(n_80), .A2(n_66), .ZN(n_18_79));
   NAND2_X1 i_18_100 (.A1(n_82), .A2(multiplicand[19]), .ZN(n_18_80));
   NAND4_X1 i_18_101 (.A1(n_18_77), .A2(n_18_78), .A3(n_18_79), .A4(n_18_80), 
      .ZN(n_103));
   NAND2_X1 i_18_102 (.A1(n_81), .A2(multiplicand[21]), .ZN(n_18_81));
   NAND2_X1 i_18_103 (.A1(n_79), .A2(n_68), .ZN(n_18_82));
   NAND2_X1 i_18_104 (.A1(n_80), .A2(n_67), .ZN(n_18_83));
   NAND2_X1 i_18_105 (.A1(n_82), .A2(multiplicand[20]), .ZN(n_18_84));
   NAND4_X1 i_18_106 (.A1(n_18_81), .A2(n_18_82), .A3(n_18_83), .A4(n_18_84), 
      .ZN(n_104));
   NAND2_X1 i_18_107 (.A1(n_81), .A2(multiplicand[22]), .ZN(n_18_85));
   NAND2_X1 i_18_108 (.A1(n_79), .A2(n_69), .ZN(n_18_86));
   NAND2_X1 i_18_109 (.A1(n_80), .A2(n_68), .ZN(n_18_87));
   NAND2_X1 i_18_110 (.A1(n_82), .A2(multiplicand[21]), .ZN(n_18_88));
   NAND4_X1 i_18_111 (.A1(n_18_85), .A2(n_18_86), .A3(n_18_87), .A4(n_18_88), 
      .ZN(n_105));
   NAND2_X1 i_18_112 (.A1(n_81), .A2(multiplicand[23]), .ZN(n_18_89));
   NAND2_X1 i_18_113 (.A1(n_79), .A2(n_70), .ZN(n_18_90));
   NAND2_X1 i_18_114 (.A1(n_80), .A2(n_69), .ZN(n_18_91));
   NAND2_X1 i_18_115 (.A1(n_82), .A2(multiplicand[22]), .ZN(n_18_92));
   NAND4_X1 i_18_116 (.A1(n_18_89), .A2(n_18_90), .A3(n_18_91), .A4(n_18_92), 
      .ZN(n_106));
   NAND2_X1 i_18_117 (.A1(n_81), .A2(multiplicand[24]), .ZN(n_18_93));
   NAND2_X1 i_18_118 (.A1(n_79), .A2(n_71), .ZN(n_18_94));
   NAND2_X1 i_18_119 (.A1(n_80), .A2(n_70), .ZN(n_18_95));
   NAND2_X1 i_18_120 (.A1(n_82), .A2(multiplicand[23]), .ZN(n_18_96));
   NAND4_X1 i_18_121 (.A1(n_18_93), .A2(n_18_94), .A3(n_18_95), .A4(n_18_96), 
      .ZN(n_107));
   NAND2_X1 i_18_122 (.A1(n_81), .A2(multiplicand[25]), .ZN(n_18_97));
   NAND2_X1 i_18_123 (.A1(n_79), .A2(n_72), .ZN(n_18_98));
   NAND2_X1 i_18_124 (.A1(n_80), .A2(n_71), .ZN(n_18_99));
   NAND2_X1 i_18_125 (.A1(n_82), .A2(multiplicand[24]), .ZN(n_18_100));
   NAND4_X1 i_18_126 (.A1(n_18_97), .A2(n_18_98), .A3(n_18_99), .A4(n_18_100), 
      .ZN(n_108));
   NAND2_X1 i_18_127 (.A1(n_81), .A2(multiplicand[26]), .ZN(n_18_101));
   NAND2_X1 i_18_128 (.A1(n_79), .A2(n_73), .ZN(n_18_102));
   NAND2_X1 i_18_129 (.A1(n_80), .A2(n_72), .ZN(n_18_103));
   NAND2_X1 i_18_130 (.A1(n_82), .A2(multiplicand[25]), .ZN(n_18_104));
   NAND4_X1 i_18_131 (.A1(n_18_101), .A2(n_18_102), .A3(n_18_103), .A4(n_18_104), 
      .ZN(n_109));
   NAND2_X1 i_18_132 (.A1(n_81), .A2(multiplicand[27]), .ZN(n_18_105));
   NAND2_X1 i_18_133 (.A1(n_79), .A2(n_74), .ZN(n_18_106));
   NAND2_X1 i_18_134 (.A1(n_80), .A2(n_73), .ZN(n_18_107));
   NAND2_X1 i_18_135 (.A1(n_82), .A2(multiplicand[26]), .ZN(n_18_108));
   NAND4_X1 i_18_136 (.A1(n_18_105), .A2(n_18_106), .A3(n_18_107), .A4(n_18_108), 
      .ZN(n_110));
   NAND2_X1 i_18_137 (.A1(n_81), .A2(multiplicand[28]), .ZN(n_18_109));
   NAND2_X1 i_18_138 (.A1(n_79), .A2(n_75), .ZN(n_18_110));
   NAND2_X1 i_18_139 (.A1(n_80), .A2(n_74), .ZN(n_18_111));
   NAND2_X1 i_18_140 (.A1(n_82), .A2(multiplicand[27]), .ZN(n_18_112));
   NAND4_X1 i_18_141 (.A1(n_18_109), .A2(n_18_110), .A3(n_18_111), .A4(n_18_112), 
      .ZN(n_111));
   NAND2_X1 i_18_142 (.A1(n_81), .A2(multiplicand[29]), .ZN(n_18_113));
   NAND2_X1 i_18_143 (.A1(n_79), .A2(n_76), .ZN(n_18_114));
   NAND2_X1 i_18_144 (.A1(n_80), .A2(n_75), .ZN(n_18_115));
   NAND2_X1 i_18_145 (.A1(n_82), .A2(multiplicand[28]), .ZN(n_18_116));
   NAND4_X1 i_18_146 (.A1(n_18_113), .A2(n_18_114), .A3(n_18_115), .A4(n_18_116), 
      .ZN(n_112));
   NAND2_X1 i_18_147 (.A1(n_81), .A2(multiplicand[30]), .ZN(n_18_117));
   NAND2_X1 i_18_148 (.A1(n_79), .A2(n_77), .ZN(n_18_118));
   NAND2_X1 i_18_149 (.A1(n_80), .A2(n_76), .ZN(n_18_119));
   NAND2_X1 i_18_150 (.A1(n_82), .A2(multiplicand[29]), .ZN(n_18_120));
   NAND4_X1 i_18_151 (.A1(n_18_117), .A2(n_18_118), .A3(n_18_119), .A4(n_18_120), 
      .ZN(n_113));
   NAND2_X1 i_18_152 (.A1(n_81), .A2(multiplicand[31]), .ZN(n_18_121));
   NAND2_X1 i_18_153 (.A1(n_79), .A2(n_78), .ZN(n_18_122));
   NAND2_X1 i_18_154 (.A1(n_80), .A2(n_77), .ZN(n_18_123));
   NAND2_X1 i_18_155 (.A1(n_82), .A2(multiplicand[30]), .ZN(n_18_124));
   NAND4_X1 i_18_156 (.A1(n_18_121), .A2(n_18_122), .A3(n_18_123), .A4(n_18_124), 
      .ZN(n_114));
   NAND2_X1 i_18_157 (.A1(n_80), .A2(n_78), .ZN(n_18_125));
   NAND2_X1 i_18_158 (.A1(n_82), .A2(multiplicand[31]), .ZN(n_18_126));
   NAND4_X1 i_18_159 (.A1(n_18_121), .A2(n_18_122), .A3(n_18_125), .A4(n_18_126), 
      .ZN(n_115));
   INV_X1 i_19_0 (.A(n_3), .ZN(n_19_0));
   AND3_X1 i_19_1 (.A1(n_19_0), .A2(n_4), .A3(n_5), .ZN(n_116));
   INV_X1 i_19_2 (.A(n_4), .ZN(n_19_1));
   AND3_X1 i_19_3 (.A1(n_19_1), .A2(n_3), .A3(n_5), .ZN(n_117));
   NOR3_X1 i_19_4 (.A1(n_19_1), .A2(n_3), .A3(n_5), .ZN(n_118));
   NOR3_X1 i_19_5 (.A1(n_19_0), .A2(n_4), .A3(n_5), .ZN(n_119));
   AOI22_X1 i_20_0 (.A1(n_118), .A2(multiplicand[0]), .B1(n_116), .B2(
      multiplicand[0]), .ZN(n_20_0));
   INV_X1 i_20_1 (.A(n_20_0), .ZN(n_120));
   NAND2_X1 i_20_2 (.A1(n_118), .A2(multiplicand[1]), .ZN(n_20_1));
   NAND2_X1 i_20_3 (.A1(n_116), .A2(n_48), .ZN(n_20_2));
   NAND2_X1 i_20_4 (.A1(n_117), .A2(multiplicand[0]), .ZN(n_20_3));
   NAND2_X1 i_20_5 (.A1(n_119), .A2(multiplicand[0]), .ZN(n_20_4));
   NAND4_X1 i_20_6 (.A1(n_20_1), .A2(n_20_2), .A3(n_20_3), .A4(n_20_4), .ZN(
      n_121));
   NAND2_X1 i_20_7 (.A1(n_118), .A2(multiplicand[2]), .ZN(n_20_5));
   NAND2_X1 i_20_8 (.A1(n_116), .A2(n_49), .ZN(n_20_6));
   NAND2_X1 i_20_9 (.A1(n_117), .A2(n_48), .ZN(n_20_7));
   NAND2_X1 i_20_10 (.A1(n_119), .A2(multiplicand[1]), .ZN(n_20_8));
   NAND4_X1 i_20_11 (.A1(n_20_5), .A2(n_20_6), .A3(n_20_7), .A4(n_20_8), 
      .ZN(n_122));
   NAND2_X1 i_20_12 (.A1(n_118), .A2(multiplicand[3]), .ZN(n_20_9));
   NAND2_X1 i_20_13 (.A1(n_116), .A2(n_50), .ZN(n_20_10));
   NAND2_X1 i_20_14 (.A1(n_117), .A2(n_49), .ZN(n_20_11));
   NAND2_X1 i_20_15 (.A1(n_119), .A2(multiplicand[2]), .ZN(n_20_12));
   NAND4_X1 i_20_16 (.A1(n_20_9), .A2(n_20_10), .A3(n_20_11), .A4(n_20_12), 
      .ZN(n_123));
   NAND2_X1 i_20_17 (.A1(n_118), .A2(multiplicand[4]), .ZN(n_20_13));
   NAND2_X1 i_20_18 (.A1(n_116), .A2(n_51), .ZN(n_20_14));
   NAND2_X1 i_20_19 (.A1(n_117), .A2(n_50), .ZN(n_20_15));
   NAND2_X1 i_20_20 (.A1(n_119), .A2(multiplicand[3]), .ZN(n_20_16));
   NAND4_X1 i_20_21 (.A1(n_20_13), .A2(n_20_14), .A3(n_20_15), .A4(n_20_16), 
      .ZN(n_124));
   NAND2_X1 i_20_22 (.A1(n_118), .A2(multiplicand[5]), .ZN(n_20_17));
   NAND2_X1 i_20_23 (.A1(n_116), .A2(n_52), .ZN(n_20_18));
   NAND2_X1 i_20_24 (.A1(n_117), .A2(n_51), .ZN(n_20_19));
   NAND2_X1 i_20_25 (.A1(n_119), .A2(multiplicand[4]), .ZN(n_20_20));
   NAND4_X1 i_20_26 (.A1(n_20_17), .A2(n_20_18), .A3(n_20_19), .A4(n_20_20), 
      .ZN(n_125));
   NAND2_X1 i_20_27 (.A1(n_118), .A2(multiplicand[6]), .ZN(n_20_21));
   NAND2_X1 i_20_28 (.A1(n_116), .A2(n_53), .ZN(n_20_22));
   NAND2_X1 i_20_29 (.A1(n_117), .A2(n_52), .ZN(n_20_23));
   NAND2_X1 i_20_30 (.A1(n_119), .A2(multiplicand[5]), .ZN(n_20_24));
   NAND4_X1 i_20_31 (.A1(n_20_21), .A2(n_20_22), .A3(n_20_23), .A4(n_20_24), 
      .ZN(n_126));
   NAND2_X1 i_20_32 (.A1(n_118), .A2(multiplicand[7]), .ZN(n_20_25));
   NAND2_X1 i_20_33 (.A1(n_116), .A2(n_54), .ZN(n_20_26));
   NAND2_X1 i_20_34 (.A1(n_117), .A2(n_53), .ZN(n_20_27));
   NAND2_X1 i_20_35 (.A1(n_119), .A2(multiplicand[6]), .ZN(n_20_28));
   NAND4_X1 i_20_36 (.A1(n_20_25), .A2(n_20_26), .A3(n_20_27), .A4(n_20_28), 
      .ZN(n_127));
   NAND2_X1 i_20_37 (.A1(n_118), .A2(multiplicand[8]), .ZN(n_20_29));
   NAND2_X1 i_20_38 (.A1(n_116), .A2(n_55), .ZN(n_20_30));
   NAND2_X1 i_20_39 (.A1(n_117), .A2(n_54), .ZN(n_20_31));
   NAND2_X1 i_20_40 (.A1(n_119), .A2(multiplicand[7]), .ZN(n_20_32));
   NAND4_X1 i_20_41 (.A1(n_20_29), .A2(n_20_30), .A3(n_20_31), .A4(n_20_32), 
      .ZN(n_128));
   NAND2_X1 i_20_42 (.A1(n_118), .A2(multiplicand[9]), .ZN(n_20_33));
   NAND2_X1 i_20_43 (.A1(n_116), .A2(n_56), .ZN(n_20_34));
   NAND2_X1 i_20_44 (.A1(n_117), .A2(n_55), .ZN(n_20_35));
   NAND2_X1 i_20_45 (.A1(n_119), .A2(multiplicand[8]), .ZN(n_20_36));
   NAND4_X1 i_20_46 (.A1(n_20_33), .A2(n_20_34), .A3(n_20_35), .A4(n_20_36), 
      .ZN(n_129));
   NAND2_X1 i_20_47 (.A1(n_118), .A2(multiplicand[10]), .ZN(n_20_37));
   NAND2_X1 i_20_48 (.A1(n_116), .A2(n_57), .ZN(n_20_38));
   NAND2_X1 i_20_49 (.A1(n_117), .A2(n_56), .ZN(n_20_39));
   NAND2_X1 i_20_50 (.A1(n_119), .A2(multiplicand[9]), .ZN(n_20_40));
   NAND4_X1 i_20_51 (.A1(n_20_37), .A2(n_20_38), .A3(n_20_39), .A4(n_20_40), 
      .ZN(n_130));
   NAND2_X1 i_20_52 (.A1(n_118), .A2(multiplicand[11]), .ZN(n_20_41));
   NAND2_X1 i_20_53 (.A1(n_116), .A2(n_58), .ZN(n_20_42));
   NAND2_X1 i_20_54 (.A1(n_117), .A2(n_57), .ZN(n_20_43));
   NAND2_X1 i_20_55 (.A1(n_119), .A2(multiplicand[10]), .ZN(n_20_44));
   NAND4_X1 i_20_56 (.A1(n_20_41), .A2(n_20_42), .A3(n_20_43), .A4(n_20_44), 
      .ZN(n_131));
   NAND2_X1 i_20_57 (.A1(n_118), .A2(multiplicand[12]), .ZN(n_20_45));
   NAND2_X1 i_20_58 (.A1(n_116), .A2(n_59), .ZN(n_20_46));
   NAND2_X1 i_20_59 (.A1(n_117), .A2(n_58), .ZN(n_20_47));
   NAND2_X1 i_20_60 (.A1(n_119), .A2(multiplicand[11]), .ZN(n_20_48));
   NAND4_X1 i_20_61 (.A1(n_20_45), .A2(n_20_46), .A3(n_20_47), .A4(n_20_48), 
      .ZN(n_132));
   NAND2_X1 i_20_62 (.A1(n_118), .A2(multiplicand[13]), .ZN(n_20_49));
   NAND2_X1 i_20_63 (.A1(n_116), .A2(n_60), .ZN(n_20_50));
   NAND2_X1 i_20_64 (.A1(n_117), .A2(n_59), .ZN(n_20_51));
   NAND2_X1 i_20_65 (.A1(n_119), .A2(multiplicand[12]), .ZN(n_20_52));
   NAND4_X1 i_20_66 (.A1(n_20_49), .A2(n_20_50), .A3(n_20_51), .A4(n_20_52), 
      .ZN(n_133));
   NAND2_X1 i_20_67 (.A1(n_118), .A2(multiplicand[14]), .ZN(n_20_53));
   NAND2_X1 i_20_68 (.A1(n_116), .A2(n_61), .ZN(n_20_54));
   NAND2_X1 i_20_69 (.A1(n_117), .A2(n_60), .ZN(n_20_55));
   NAND2_X1 i_20_70 (.A1(n_119), .A2(multiplicand[13]), .ZN(n_20_56));
   NAND4_X1 i_20_71 (.A1(n_20_53), .A2(n_20_54), .A3(n_20_55), .A4(n_20_56), 
      .ZN(n_134));
   NAND2_X1 i_20_72 (.A1(n_118), .A2(multiplicand[15]), .ZN(n_20_57));
   NAND2_X1 i_20_73 (.A1(n_116), .A2(n_62), .ZN(n_20_58));
   NAND2_X1 i_20_74 (.A1(n_117), .A2(n_61), .ZN(n_20_59));
   NAND2_X1 i_20_75 (.A1(n_119), .A2(multiplicand[14]), .ZN(n_20_60));
   NAND4_X1 i_20_76 (.A1(n_20_57), .A2(n_20_58), .A3(n_20_59), .A4(n_20_60), 
      .ZN(n_135));
   NAND2_X1 i_20_77 (.A1(n_118), .A2(multiplicand[16]), .ZN(n_20_61));
   NAND2_X1 i_20_78 (.A1(n_116), .A2(n_63), .ZN(n_20_62));
   NAND2_X1 i_20_79 (.A1(n_117), .A2(n_62), .ZN(n_20_63));
   NAND2_X1 i_20_80 (.A1(n_119), .A2(multiplicand[15]), .ZN(n_20_64));
   NAND4_X1 i_20_81 (.A1(n_20_61), .A2(n_20_62), .A3(n_20_63), .A4(n_20_64), 
      .ZN(n_136));
   NAND2_X1 i_20_82 (.A1(n_118), .A2(multiplicand[17]), .ZN(n_20_65));
   NAND2_X1 i_20_83 (.A1(n_116), .A2(n_64), .ZN(n_20_66));
   NAND2_X1 i_20_84 (.A1(n_117), .A2(n_63), .ZN(n_20_67));
   NAND2_X1 i_20_85 (.A1(n_119), .A2(multiplicand[16]), .ZN(n_20_68));
   NAND4_X1 i_20_86 (.A1(n_20_65), .A2(n_20_66), .A3(n_20_67), .A4(n_20_68), 
      .ZN(n_137));
   NAND2_X1 i_20_87 (.A1(n_118), .A2(multiplicand[18]), .ZN(n_20_69));
   NAND2_X1 i_20_88 (.A1(n_116), .A2(n_65), .ZN(n_20_70));
   NAND2_X1 i_20_89 (.A1(n_117), .A2(n_64), .ZN(n_20_71));
   NAND2_X1 i_20_90 (.A1(n_119), .A2(multiplicand[17]), .ZN(n_20_72));
   NAND4_X1 i_20_91 (.A1(n_20_69), .A2(n_20_70), .A3(n_20_71), .A4(n_20_72), 
      .ZN(n_138));
   NAND2_X1 i_20_92 (.A1(n_118), .A2(multiplicand[19]), .ZN(n_20_73));
   NAND2_X1 i_20_93 (.A1(n_116), .A2(n_66), .ZN(n_20_74));
   NAND2_X1 i_20_94 (.A1(n_117), .A2(n_65), .ZN(n_20_75));
   NAND2_X1 i_20_95 (.A1(n_119), .A2(multiplicand[18]), .ZN(n_20_76));
   NAND4_X1 i_20_96 (.A1(n_20_73), .A2(n_20_74), .A3(n_20_75), .A4(n_20_76), 
      .ZN(n_139));
   NAND2_X1 i_20_97 (.A1(n_118), .A2(multiplicand[20]), .ZN(n_20_77));
   NAND2_X1 i_20_98 (.A1(n_116), .A2(n_67), .ZN(n_20_78));
   NAND2_X1 i_20_99 (.A1(n_117), .A2(n_66), .ZN(n_20_79));
   NAND2_X1 i_20_100 (.A1(n_119), .A2(multiplicand[19]), .ZN(n_20_80));
   NAND4_X1 i_20_101 (.A1(n_20_77), .A2(n_20_78), .A3(n_20_79), .A4(n_20_80), 
      .ZN(n_140));
   NAND2_X1 i_20_102 (.A1(n_118), .A2(multiplicand[21]), .ZN(n_20_81));
   NAND2_X1 i_20_103 (.A1(n_116), .A2(n_68), .ZN(n_20_82));
   NAND2_X1 i_20_104 (.A1(n_117), .A2(n_67), .ZN(n_20_83));
   NAND2_X1 i_20_105 (.A1(n_119), .A2(multiplicand[20]), .ZN(n_20_84));
   NAND4_X1 i_20_106 (.A1(n_20_81), .A2(n_20_82), .A3(n_20_83), .A4(n_20_84), 
      .ZN(n_141));
   NAND2_X1 i_20_107 (.A1(n_118), .A2(multiplicand[22]), .ZN(n_20_85));
   NAND2_X1 i_20_108 (.A1(n_116), .A2(n_69), .ZN(n_20_86));
   NAND2_X1 i_20_109 (.A1(n_117), .A2(n_68), .ZN(n_20_87));
   NAND2_X1 i_20_110 (.A1(n_119), .A2(multiplicand[21]), .ZN(n_20_88));
   NAND4_X1 i_20_111 (.A1(n_20_85), .A2(n_20_86), .A3(n_20_87), .A4(n_20_88), 
      .ZN(n_142));
   NAND2_X1 i_20_112 (.A1(n_118), .A2(multiplicand[23]), .ZN(n_20_89));
   NAND2_X1 i_20_113 (.A1(n_116), .A2(n_70), .ZN(n_20_90));
   NAND2_X1 i_20_114 (.A1(n_117), .A2(n_69), .ZN(n_20_91));
   NAND2_X1 i_20_115 (.A1(n_119), .A2(multiplicand[22]), .ZN(n_20_92));
   NAND4_X1 i_20_116 (.A1(n_20_89), .A2(n_20_90), .A3(n_20_91), .A4(n_20_92), 
      .ZN(n_143));
   NAND2_X1 i_20_117 (.A1(n_118), .A2(multiplicand[24]), .ZN(n_20_93));
   NAND2_X1 i_20_118 (.A1(n_116), .A2(n_71), .ZN(n_20_94));
   NAND2_X1 i_20_119 (.A1(n_117), .A2(n_70), .ZN(n_20_95));
   NAND2_X1 i_20_120 (.A1(n_119), .A2(multiplicand[23]), .ZN(n_20_96));
   NAND4_X1 i_20_121 (.A1(n_20_93), .A2(n_20_94), .A3(n_20_95), .A4(n_20_96), 
      .ZN(n_144));
   NAND2_X1 i_20_122 (.A1(n_118), .A2(multiplicand[25]), .ZN(n_20_97));
   NAND2_X1 i_20_123 (.A1(n_116), .A2(n_72), .ZN(n_20_98));
   NAND2_X1 i_20_124 (.A1(n_117), .A2(n_71), .ZN(n_20_99));
   NAND2_X1 i_20_125 (.A1(n_119), .A2(multiplicand[24]), .ZN(n_20_100));
   NAND4_X1 i_20_126 (.A1(n_20_97), .A2(n_20_98), .A3(n_20_99), .A4(n_20_100), 
      .ZN(n_145));
   NAND2_X1 i_20_127 (.A1(n_118), .A2(multiplicand[26]), .ZN(n_20_101));
   NAND2_X1 i_20_128 (.A1(n_116), .A2(n_73), .ZN(n_20_102));
   NAND2_X1 i_20_129 (.A1(n_117), .A2(n_72), .ZN(n_20_103));
   NAND2_X1 i_20_130 (.A1(n_119), .A2(multiplicand[25]), .ZN(n_20_104));
   NAND4_X1 i_20_131 (.A1(n_20_101), .A2(n_20_102), .A3(n_20_103), .A4(n_20_104), 
      .ZN(n_146));
   NAND2_X1 i_20_132 (.A1(n_118), .A2(multiplicand[27]), .ZN(n_20_105));
   NAND2_X1 i_20_133 (.A1(n_116), .A2(n_74), .ZN(n_20_106));
   NAND2_X1 i_20_134 (.A1(n_117), .A2(n_73), .ZN(n_20_107));
   NAND2_X1 i_20_135 (.A1(n_119), .A2(multiplicand[26]), .ZN(n_20_108));
   NAND4_X1 i_20_136 (.A1(n_20_105), .A2(n_20_106), .A3(n_20_107), .A4(n_20_108), 
      .ZN(n_147));
   NAND2_X1 i_20_137 (.A1(n_118), .A2(multiplicand[28]), .ZN(n_20_109));
   NAND2_X1 i_20_138 (.A1(n_116), .A2(n_75), .ZN(n_20_110));
   NAND2_X1 i_20_139 (.A1(n_117), .A2(n_74), .ZN(n_20_111));
   NAND2_X1 i_20_140 (.A1(n_119), .A2(multiplicand[27]), .ZN(n_20_112));
   NAND4_X1 i_20_141 (.A1(n_20_109), .A2(n_20_110), .A3(n_20_111), .A4(n_20_112), 
      .ZN(n_148));
   NAND2_X1 i_20_142 (.A1(n_118), .A2(multiplicand[29]), .ZN(n_20_113));
   NAND2_X1 i_20_143 (.A1(n_116), .A2(n_76), .ZN(n_20_114));
   NAND2_X1 i_20_144 (.A1(n_117), .A2(n_75), .ZN(n_20_115));
   NAND2_X1 i_20_145 (.A1(n_119), .A2(multiplicand[28]), .ZN(n_20_116));
   NAND4_X1 i_20_146 (.A1(n_20_113), .A2(n_20_114), .A3(n_20_115), .A4(n_20_116), 
      .ZN(n_149));
   NAND2_X1 i_20_147 (.A1(n_118), .A2(multiplicand[30]), .ZN(n_20_117));
   NAND2_X1 i_20_148 (.A1(n_116), .A2(n_77), .ZN(n_20_118));
   NAND2_X1 i_20_149 (.A1(n_117), .A2(n_76), .ZN(n_20_119));
   NAND2_X1 i_20_150 (.A1(n_119), .A2(multiplicand[29]), .ZN(n_20_120));
   NAND4_X1 i_20_151 (.A1(n_20_117), .A2(n_20_118), .A3(n_20_119), .A4(n_20_120), 
      .ZN(n_150));
   NAND2_X1 i_20_152 (.A1(n_118), .A2(multiplicand[31]), .ZN(n_20_121));
   NAND2_X1 i_20_153 (.A1(n_116), .A2(n_78), .ZN(n_20_122));
   NAND2_X1 i_20_154 (.A1(n_117), .A2(n_77), .ZN(n_20_123));
   NAND2_X1 i_20_155 (.A1(n_119), .A2(multiplicand[30]), .ZN(n_20_124));
   NAND4_X1 i_20_156 (.A1(n_20_121), .A2(n_20_122), .A3(n_20_123), .A4(n_20_124), 
      .ZN(n_151));
   NAND2_X1 i_20_157 (.A1(n_117), .A2(n_78), .ZN(n_20_125));
   NAND2_X1 i_20_158 (.A1(n_119), .A2(multiplicand[31]), .ZN(n_20_126));
   NAND4_X1 i_20_159 (.A1(n_20_121), .A2(n_20_122), .A3(n_20_125), .A4(n_20_126), 
      .ZN(n_152));
   INV_X1 i_21_0 (.A(n_6), .ZN(n_21_0));
   AND3_X1 i_21_1 (.A1(n_21_0), .A2(n_7), .A3(n_8), .ZN(n_153));
   INV_X1 i_21_2 (.A(n_7), .ZN(n_21_1));
   AND3_X1 i_21_3 (.A1(n_21_1), .A2(n_6), .A3(n_8), .ZN(n_154));
   NOR3_X1 i_21_4 (.A1(n_21_1), .A2(n_6), .A3(n_8), .ZN(n_155));
   NOR3_X1 i_21_5 (.A1(n_21_0), .A2(n_7), .A3(n_8), .ZN(n_156));
   AOI22_X1 i_22_0 (.A1(n_155), .A2(multiplicand[0]), .B1(n_153), .B2(
      multiplicand[0]), .ZN(n_22_0));
   INV_X1 i_22_1 (.A(n_22_0), .ZN(n_157));
   NAND2_X1 i_22_2 (.A1(n_155), .A2(multiplicand[1]), .ZN(n_22_1));
   NAND2_X1 i_22_3 (.A1(n_153), .A2(n_48), .ZN(n_22_2));
   NAND2_X1 i_22_4 (.A1(n_154), .A2(multiplicand[0]), .ZN(n_22_3));
   NAND2_X1 i_22_5 (.A1(n_156), .A2(multiplicand[0]), .ZN(n_22_4));
   NAND4_X1 i_22_6 (.A1(n_22_1), .A2(n_22_2), .A3(n_22_3), .A4(n_22_4), .ZN(
      n_158));
   NAND2_X1 i_22_7 (.A1(n_155), .A2(multiplicand[2]), .ZN(n_22_5));
   NAND2_X1 i_22_8 (.A1(n_153), .A2(n_49), .ZN(n_22_6));
   NAND2_X1 i_22_9 (.A1(n_154), .A2(n_48), .ZN(n_22_7));
   NAND2_X1 i_22_10 (.A1(n_156), .A2(multiplicand[1]), .ZN(n_22_8));
   NAND4_X1 i_22_11 (.A1(n_22_5), .A2(n_22_6), .A3(n_22_7), .A4(n_22_8), 
      .ZN(n_159));
   NAND2_X1 i_22_12 (.A1(n_155), .A2(multiplicand[3]), .ZN(n_22_9));
   NAND2_X1 i_22_13 (.A1(n_153), .A2(n_50), .ZN(n_22_10));
   NAND2_X1 i_22_14 (.A1(n_154), .A2(n_49), .ZN(n_22_11));
   NAND2_X1 i_22_15 (.A1(n_156), .A2(multiplicand[2]), .ZN(n_22_12));
   NAND4_X1 i_22_16 (.A1(n_22_9), .A2(n_22_10), .A3(n_22_11), .A4(n_22_12), 
      .ZN(n_160));
   NAND2_X1 i_22_17 (.A1(n_155), .A2(multiplicand[4]), .ZN(n_22_13));
   NAND2_X1 i_22_18 (.A1(n_153), .A2(n_51), .ZN(n_22_14));
   NAND2_X1 i_22_19 (.A1(n_154), .A2(n_50), .ZN(n_22_15));
   NAND2_X1 i_22_20 (.A1(n_156), .A2(multiplicand[3]), .ZN(n_22_16));
   NAND4_X1 i_22_21 (.A1(n_22_13), .A2(n_22_14), .A3(n_22_15), .A4(n_22_16), 
      .ZN(n_161));
   NAND2_X1 i_22_22 (.A1(n_155), .A2(multiplicand[5]), .ZN(n_22_17));
   NAND2_X1 i_22_23 (.A1(n_153), .A2(n_52), .ZN(n_22_18));
   NAND2_X1 i_22_24 (.A1(n_154), .A2(n_51), .ZN(n_22_19));
   NAND2_X1 i_22_25 (.A1(n_156), .A2(multiplicand[4]), .ZN(n_22_20));
   NAND4_X1 i_22_26 (.A1(n_22_17), .A2(n_22_18), .A3(n_22_19), .A4(n_22_20), 
      .ZN(n_162));
   NAND2_X1 i_22_27 (.A1(n_155), .A2(multiplicand[6]), .ZN(n_22_21));
   NAND2_X1 i_22_28 (.A1(n_153), .A2(n_53), .ZN(n_22_22));
   NAND2_X1 i_22_29 (.A1(n_154), .A2(n_52), .ZN(n_22_23));
   NAND2_X1 i_22_30 (.A1(n_156), .A2(multiplicand[5]), .ZN(n_22_24));
   NAND4_X1 i_22_31 (.A1(n_22_21), .A2(n_22_22), .A3(n_22_23), .A4(n_22_24), 
      .ZN(n_163));
   NAND2_X1 i_22_32 (.A1(n_155), .A2(multiplicand[7]), .ZN(n_22_25));
   NAND2_X1 i_22_33 (.A1(n_153), .A2(n_54), .ZN(n_22_26));
   NAND2_X1 i_22_34 (.A1(n_154), .A2(n_53), .ZN(n_22_27));
   NAND2_X1 i_22_35 (.A1(n_156), .A2(multiplicand[6]), .ZN(n_22_28));
   NAND4_X1 i_22_36 (.A1(n_22_25), .A2(n_22_26), .A3(n_22_27), .A4(n_22_28), 
      .ZN(n_164));
   NAND2_X1 i_22_37 (.A1(n_155), .A2(multiplicand[8]), .ZN(n_22_29));
   NAND2_X1 i_22_38 (.A1(n_153), .A2(n_55), .ZN(n_22_30));
   NAND2_X1 i_22_39 (.A1(n_154), .A2(n_54), .ZN(n_22_31));
   NAND2_X1 i_22_40 (.A1(n_156), .A2(multiplicand[7]), .ZN(n_22_32));
   NAND4_X1 i_22_41 (.A1(n_22_29), .A2(n_22_30), .A3(n_22_31), .A4(n_22_32), 
      .ZN(n_165));
   NAND2_X1 i_22_42 (.A1(n_155), .A2(multiplicand[9]), .ZN(n_22_33));
   NAND2_X1 i_22_43 (.A1(n_153), .A2(n_56), .ZN(n_22_34));
   NAND2_X1 i_22_44 (.A1(n_154), .A2(n_55), .ZN(n_22_35));
   NAND2_X1 i_22_45 (.A1(n_156), .A2(multiplicand[8]), .ZN(n_22_36));
   NAND4_X1 i_22_46 (.A1(n_22_33), .A2(n_22_34), .A3(n_22_35), .A4(n_22_36), 
      .ZN(n_166));
   NAND2_X1 i_22_47 (.A1(n_155), .A2(multiplicand[10]), .ZN(n_22_37));
   NAND2_X1 i_22_48 (.A1(n_153), .A2(n_57), .ZN(n_22_38));
   NAND2_X1 i_22_49 (.A1(n_154), .A2(n_56), .ZN(n_22_39));
   NAND2_X1 i_22_50 (.A1(n_156), .A2(multiplicand[9]), .ZN(n_22_40));
   NAND4_X1 i_22_51 (.A1(n_22_37), .A2(n_22_38), .A3(n_22_39), .A4(n_22_40), 
      .ZN(n_167));
   NAND2_X1 i_22_52 (.A1(n_155), .A2(multiplicand[11]), .ZN(n_22_41));
   NAND2_X1 i_22_53 (.A1(n_153), .A2(n_58), .ZN(n_22_42));
   NAND2_X1 i_22_54 (.A1(n_154), .A2(n_57), .ZN(n_22_43));
   NAND2_X1 i_22_55 (.A1(n_156), .A2(multiplicand[10]), .ZN(n_22_44));
   NAND4_X1 i_22_56 (.A1(n_22_41), .A2(n_22_42), .A3(n_22_43), .A4(n_22_44), 
      .ZN(n_168));
   NAND2_X1 i_22_57 (.A1(n_155), .A2(multiplicand[12]), .ZN(n_22_45));
   NAND2_X1 i_22_58 (.A1(n_153), .A2(n_59), .ZN(n_22_46));
   NAND2_X1 i_22_59 (.A1(n_154), .A2(n_58), .ZN(n_22_47));
   NAND2_X1 i_22_60 (.A1(n_156), .A2(multiplicand[11]), .ZN(n_22_48));
   NAND4_X1 i_22_61 (.A1(n_22_45), .A2(n_22_46), .A3(n_22_47), .A4(n_22_48), 
      .ZN(n_169));
   NAND2_X1 i_22_62 (.A1(n_155), .A2(multiplicand[13]), .ZN(n_22_49));
   NAND2_X1 i_22_63 (.A1(n_153), .A2(n_60), .ZN(n_22_50));
   NAND2_X1 i_22_64 (.A1(n_154), .A2(n_59), .ZN(n_22_51));
   NAND2_X1 i_22_65 (.A1(n_156), .A2(multiplicand[12]), .ZN(n_22_52));
   NAND4_X1 i_22_66 (.A1(n_22_49), .A2(n_22_50), .A3(n_22_51), .A4(n_22_52), 
      .ZN(n_170));
   NAND2_X1 i_22_67 (.A1(n_155), .A2(multiplicand[14]), .ZN(n_22_53));
   NAND2_X1 i_22_68 (.A1(n_153), .A2(n_61), .ZN(n_22_54));
   NAND2_X1 i_22_69 (.A1(n_154), .A2(n_60), .ZN(n_22_55));
   NAND2_X1 i_22_70 (.A1(n_156), .A2(multiplicand[13]), .ZN(n_22_56));
   NAND4_X1 i_22_71 (.A1(n_22_53), .A2(n_22_54), .A3(n_22_55), .A4(n_22_56), 
      .ZN(n_171));
   NAND2_X1 i_22_72 (.A1(n_155), .A2(multiplicand[15]), .ZN(n_22_57));
   NAND2_X1 i_22_73 (.A1(n_153), .A2(n_62), .ZN(n_22_58));
   NAND2_X1 i_22_74 (.A1(n_154), .A2(n_61), .ZN(n_22_59));
   NAND2_X1 i_22_75 (.A1(n_156), .A2(multiplicand[14]), .ZN(n_22_60));
   NAND4_X1 i_22_76 (.A1(n_22_57), .A2(n_22_58), .A3(n_22_59), .A4(n_22_60), 
      .ZN(n_172));
   NAND2_X1 i_22_77 (.A1(n_155), .A2(multiplicand[16]), .ZN(n_22_61));
   NAND2_X1 i_22_78 (.A1(n_153), .A2(n_63), .ZN(n_22_62));
   NAND2_X1 i_22_79 (.A1(n_154), .A2(n_62), .ZN(n_22_63));
   NAND2_X1 i_22_80 (.A1(n_156), .A2(multiplicand[15]), .ZN(n_22_64));
   NAND4_X1 i_22_81 (.A1(n_22_61), .A2(n_22_62), .A3(n_22_63), .A4(n_22_64), 
      .ZN(n_173));
   NAND2_X1 i_22_82 (.A1(n_155), .A2(multiplicand[17]), .ZN(n_22_65));
   NAND2_X1 i_22_83 (.A1(n_153), .A2(n_64), .ZN(n_22_66));
   NAND2_X1 i_22_84 (.A1(n_154), .A2(n_63), .ZN(n_22_67));
   NAND2_X1 i_22_85 (.A1(n_156), .A2(multiplicand[16]), .ZN(n_22_68));
   NAND4_X1 i_22_86 (.A1(n_22_65), .A2(n_22_66), .A3(n_22_67), .A4(n_22_68), 
      .ZN(n_174));
   NAND2_X1 i_22_87 (.A1(n_155), .A2(multiplicand[18]), .ZN(n_22_69));
   NAND2_X1 i_22_88 (.A1(n_153), .A2(n_65), .ZN(n_22_70));
   NAND2_X1 i_22_89 (.A1(n_154), .A2(n_64), .ZN(n_22_71));
   NAND2_X1 i_22_90 (.A1(n_156), .A2(multiplicand[17]), .ZN(n_22_72));
   NAND4_X1 i_22_91 (.A1(n_22_69), .A2(n_22_70), .A3(n_22_71), .A4(n_22_72), 
      .ZN(n_175));
   NAND2_X1 i_22_92 (.A1(n_155), .A2(multiplicand[19]), .ZN(n_22_73));
   NAND2_X1 i_22_93 (.A1(n_153), .A2(n_66), .ZN(n_22_74));
   NAND2_X1 i_22_94 (.A1(n_154), .A2(n_65), .ZN(n_22_75));
   NAND2_X1 i_22_95 (.A1(n_156), .A2(multiplicand[18]), .ZN(n_22_76));
   NAND4_X1 i_22_96 (.A1(n_22_73), .A2(n_22_74), .A3(n_22_75), .A4(n_22_76), 
      .ZN(n_176));
   NAND2_X1 i_22_97 (.A1(n_155), .A2(multiplicand[20]), .ZN(n_22_77));
   NAND2_X1 i_22_98 (.A1(n_153), .A2(n_67), .ZN(n_22_78));
   NAND2_X1 i_22_99 (.A1(n_154), .A2(n_66), .ZN(n_22_79));
   NAND2_X1 i_22_100 (.A1(n_156), .A2(multiplicand[19]), .ZN(n_22_80));
   NAND4_X1 i_22_101 (.A1(n_22_77), .A2(n_22_78), .A3(n_22_79), .A4(n_22_80), 
      .ZN(n_177));
   NAND2_X1 i_22_102 (.A1(n_155), .A2(multiplicand[21]), .ZN(n_22_81));
   NAND2_X1 i_22_103 (.A1(n_153), .A2(n_68), .ZN(n_22_82));
   NAND2_X1 i_22_104 (.A1(n_154), .A2(n_67), .ZN(n_22_83));
   NAND2_X1 i_22_105 (.A1(n_156), .A2(multiplicand[20]), .ZN(n_22_84));
   NAND4_X1 i_22_106 (.A1(n_22_81), .A2(n_22_82), .A3(n_22_83), .A4(n_22_84), 
      .ZN(n_178));
   NAND2_X1 i_22_107 (.A1(n_155), .A2(multiplicand[22]), .ZN(n_22_85));
   NAND2_X1 i_22_108 (.A1(n_153), .A2(n_69), .ZN(n_22_86));
   NAND2_X1 i_22_109 (.A1(n_154), .A2(n_68), .ZN(n_22_87));
   NAND2_X1 i_22_110 (.A1(n_156), .A2(multiplicand[21]), .ZN(n_22_88));
   NAND4_X1 i_22_111 (.A1(n_22_85), .A2(n_22_86), .A3(n_22_87), .A4(n_22_88), 
      .ZN(n_179));
   NAND2_X1 i_22_112 (.A1(n_155), .A2(multiplicand[23]), .ZN(n_22_89));
   NAND2_X1 i_22_113 (.A1(n_153), .A2(n_70), .ZN(n_22_90));
   NAND2_X1 i_22_114 (.A1(n_154), .A2(n_69), .ZN(n_22_91));
   NAND2_X1 i_22_115 (.A1(n_156), .A2(multiplicand[22]), .ZN(n_22_92));
   NAND4_X1 i_22_116 (.A1(n_22_89), .A2(n_22_90), .A3(n_22_91), .A4(n_22_92), 
      .ZN(n_180));
   NAND2_X1 i_22_117 (.A1(n_155), .A2(multiplicand[24]), .ZN(n_22_93));
   NAND2_X1 i_22_118 (.A1(n_153), .A2(n_71), .ZN(n_22_94));
   NAND2_X1 i_22_119 (.A1(n_154), .A2(n_70), .ZN(n_22_95));
   NAND2_X1 i_22_120 (.A1(n_156), .A2(multiplicand[23]), .ZN(n_22_96));
   NAND4_X1 i_22_121 (.A1(n_22_93), .A2(n_22_94), .A3(n_22_95), .A4(n_22_96), 
      .ZN(n_181));
   NAND2_X1 i_22_122 (.A1(n_155), .A2(multiplicand[25]), .ZN(n_22_97));
   NAND2_X1 i_22_123 (.A1(n_153), .A2(n_72), .ZN(n_22_98));
   NAND2_X1 i_22_124 (.A1(n_154), .A2(n_71), .ZN(n_22_99));
   NAND2_X1 i_22_125 (.A1(n_156), .A2(multiplicand[24]), .ZN(n_22_100));
   NAND4_X1 i_22_126 (.A1(n_22_97), .A2(n_22_98), .A3(n_22_99), .A4(n_22_100), 
      .ZN(n_182));
   NAND2_X1 i_22_127 (.A1(n_155), .A2(multiplicand[26]), .ZN(n_22_101));
   NAND2_X1 i_22_128 (.A1(n_153), .A2(n_73), .ZN(n_22_102));
   NAND2_X1 i_22_129 (.A1(n_154), .A2(n_72), .ZN(n_22_103));
   NAND2_X1 i_22_130 (.A1(n_156), .A2(multiplicand[25]), .ZN(n_22_104));
   NAND4_X1 i_22_131 (.A1(n_22_101), .A2(n_22_102), .A3(n_22_103), .A4(n_22_104), 
      .ZN(n_183));
   NAND2_X1 i_22_132 (.A1(n_155), .A2(multiplicand[27]), .ZN(n_22_105));
   NAND2_X1 i_22_133 (.A1(n_153), .A2(n_74), .ZN(n_22_106));
   NAND2_X1 i_22_134 (.A1(n_154), .A2(n_73), .ZN(n_22_107));
   NAND2_X1 i_22_135 (.A1(n_156), .A2(multiplicand[26]), .ZN(n_22_108));
   NAND4_X1 i_22_136 (.A1(n_22_105), .A2(n_22_106), .A3(n_22_107), .A4(n_22_108), 
      .ZN(n_184));
   NAND2_X1 i_22_137 (.A1(n_155), .A2(multiplicand[28]), .ZN(n_22_109));
   NAND2_X1 i_22_138 (.A1(n_153), .A2(n_75), .ZN(n_22_110));
   NAND2_X1 i_22_139 (.A1(n_154), .A2(n_74), .ZN(n_22_111));
   NAND2_X1 i_22_140 (.A1(n_156), .A2(multiplicand[27]), .ZN(n_22_112));
   NAND4_X1 i_22_141 (.A1(n_22_109), .A2(n_22_110), .A3(n_22_111), .A4(n_22_112), 
      .ZN(n_185));
   NAND2_X1 i_22_142 (.A1(n_155), .A2(multiplicand[29]), .ZN(n_22_113));
   NAND2_X1 i_22_143 (.A1(n_153), .A2(n_76), .ZN(n_22_114));
   NAND2_X1 i_22_144 (.A1(n_154), .A2(n_75), .ZN(n_22_115));
   NAND2_X1 i_22_145 (.A1(n_156), .A2(multiplicand[28]), .ZN(n_22_116));
   NAND4_X1 i_22_146 (.A1(n_22_113), .A2(n_22_114), .A3(n_22_115), .A4(n_22_116), 
      .ZN(n_186));
   NAND2_X1 i_22_147 (.A1(n_155), .A2(multiplicand[30]), .ZN(n_22_117));
   NAND2_X1 i_22_148 (.A1(n_153), .A2(n_77), .ZN(n_22_118));
   NAND2_X1 i_22_149 (.A1(n_154), .A2(n_76), .ZN(n_22_119));
   NAND2_X1 i_22_150 (.A1(n_156), .A2(multiplicand[29]), .ZN(n_22_120));
   NAND4_X1 i_22_151 (.A1(n_22_117), .A2(n_22_118), .A3(n_22_119), .A4(n_22_120), 
      .ZN(n_187));
   NAND2_X1 i_22_152 (.A1(n_155), .A2(multiplicand[31]), .ZN(n_22_121));
   NAND2_X1 i_22_153 (.A1(n_153), .A2(n_78), .ZN(n_22_122));
   NAND2_X1 i_22_154 (.A1(n_154), .A2(n_77), .ZN(n_22_123));
   NAND2_X1 i_22_155 (.A1(n_156), .A2(multiplicand[30]), .ZN(n_22_124));
   NAND4_X1 i_22_156 (.A1(n_22_121), .A2(n_22_122), .A3(n_22_123), .A4(n_22_124), 
      .ZN(n_188));
   NAND2_X1 i_22_157 (.A1(n_154), .A2(n_78), .ZN(n_22_125));
   NAND2_X1 i_22_158 (.A1(n_156), .A2(multiplicand[31]), .ZN(n_22_126));
   NAND4_X1 i_22_159 (.A1(n_22_121), .A2(n_22_122), .A3(n_22_125), .A4(n_22_126), 
      .ZN(n_189));
   INV_X1 i_23_0 (.A(n_9), .ZN(n_23_0));
   AND3_X1 i_23_1 (.A1(n_23_0), .A2(n_10), .A3(n_11), .ZN(n_190));
   INV_X1 i_23_2 (.A(n_10), .ZN(n_23_1));
   AND3_X1 i_23_3 (.A1(n_23_1), .A2(n_9), .A3(n_11), .ZN(n_191));
   NOR3_X1 i_23_4 (.A1(n_23_1), .A2(n_9), .A3(n_11), .ZN(n_192));
   NOR3_X1 i_23_5 (.A1(n_23_0), .A2(n_10), .A3(n_11), .ZN(n_193));
   AOI22_X1 i_24_0 (.A1(n_192), .A2(multiplicand[0]), .B1(n_190), .B2(
      multiplicand[0]), .ZN(n_24_0));
   INV_X1 i_24_1 (.A(n_24_0), .ZN(n_194));
   NAND2_X1 i_24_2 (.A1(n_192), .A2(multiplicand[1]), .ZN(n_24_1));
   NAND2_X1 i_24_3 (.A1(n_190), .A2(n_48), .ZN(n_24_2));
   NAND2_X1 i_24_4 (.A1(n_191), .A2(multiplicand[0]), .ZN(n_24_3));
   NAND2_X1 i_24_5 (.A1(n_193), .A2(multiplicand[0]), .ZN(n_24_4));
   NAND4_X1 i_24_6 (.A1(n_24_1), .A2(n_24_2), .A3(n_24_3), .A4(n_24_4), .ZN(
      n_195));
   NAND2_X1 i_24_7 (.A1(n_192), .A2(multiplicand[2]), .ZN(n_24_5));
   NAND2_X1 i_24_8 (.A1(n_190), .A2(n_49), .ZN(n_24_6));
   NAND2_X1 i_24_9 (.A1(n_191), .A2(n_48), .ZN(n_24_7));
   NAND2_X1 i_24_10 (.A1(n_193), .A2(multiplicand[1]), .ZN(n_24_8));
   NAND4_X1 i_24_11 (.A1(n_24_5), .A2(n_24_6), .A3(n_24_7), .A4(n_24_8), 
      .ZN(n_196));
   NAND2_X1 i_24_12 (.A1(n_192), .A2(multiplicand[3]), .ZN(n_24_9));
   NAND2_X1 i_24_13 (.A1(n_190), .A2(n_50), .ZN(n_24_10));
   NAND2_X1 i_24_14 (.A1(n_191), .A2(n_49), .ZN(n_24_11));
   NAND2_X1 i_24_15 (.A1(n_193), .A2(multiplicand[2]), .ZN(n_24_12));
   NAND4_X1 i_24_16 (.A1(n_24_9), .A2(n_24_10), .A3(n_24_11), .A4(n_24_12), 
      .ZN(n_197));
   NAND2_X1 i_24_17 (.A1(n_192), .A2(multiplicand[4]), .ZN(n_24_13));
   NAND2_X1 i_24_18 (.A1(n_190), .A2(n_51), .ZN(n_24_14));
   NAND2_X1 i_24_19 (.A1(n_191), .A2(n_50), .ZN(n_24_15));
   NAND2_X1 i_24_20 (.A1(n_193), .A2(multiplicand[3]), .ZN(n_24_16));
   NAND4_X1 i_24_21 (.A1(n_24_13), .A2(n_24_14), .A3(n_24_15), .A4(n_24_16), 
      .ZN(n_198));
   NAND2_X1 i_24_22 (.A1(n_192), .A2(multiplicand[5]), .ZN(n_24_17));
   NAND2_X1 i_24_23 (.A1(n_190), .A2(n_52), .ZN(n_24_18));
   NAND2_X1 i_24_24 (.A1(n_191), .A2(n_51), .ZN(n_24_19));
   NAND2_X1 i_24_25 (.A1(n_193), .A2(multiplicand[4]), .ZN(n_24_20));
   NAND4_X1 i_24_26 (.A1(n_24_17), .A2(n_24_18), .A3(n_24_19), .A4(n_24_20), 
      .ZN(n_199));
   NAND2_X1 i_24_27 (.A1(n_192), .A2(multiplicand[6]), .ZN(n_24_21));
   NAND2_X1 i_24_28 (.A1(n_190), .A2(n_53), .ZN(n_24_22));
   NAND2_X1 i_24_29 (.A1(n_191), .A2(n_52), .ZN(n_24_23));
   NAND2_X1 i_24_30 (.A1(n_193), .A2(multiplicand[5]), .ZN(n_24_24));
   NAND4_X1 i_24_31 (.A1(n_24_21), .A2(n_24_22), .A3(n_24_23), .A4(n_24_24), 
      .ZN(n_200));
   NAND2_X1 i_24_32 (.A1(n_192), .A2(multiplicand[7]), .ZN(n_24_25));
   NAND2_X1 i_24_33 (.A1(n_190), .A2(n_54), .ZN(n_24_26));
   NAND2_X1 i_24_34 (.A1(n_191), .A2(n_53), .ZN(n_24_27));
   NAND2_X1 i_24_35 (.A1(n_193), .A2(multiplicand[6]), .ZN(n_24_28));
   NAND4_X1 i_24_36 (.A1(n_24_25), .A2(n_24_26), .A3(n_24_27), .A4(n_24_28), 
      .ZN(n_201));
   NAND2_X1 i_24_37 (.A1(n_192), .A2(multiplicand[8]), .ZN(n_24_29));
   NAND2_X1 i_24_38 (.A1(n_190), .A2(n_55), .ZN(n_24_30));
   NAND2_X1 i_24_39 (.A1(n_191), .A2(n_54), .ZN(n_24_31));
   NAND2_X1 i_24_40 (.A1(n_193), .A2(multiplicand[7]), .ZN(n_24_32));
   NAND4_X1 i_24_41 (.A1(n_24_29), .A2(n_24_30), .A3(n_24_31), .A4(n_24_32), 
      .ZN(n_202));
   NAND2_X1 i_24_42 (.A1(n_192), .A2(multiplicand[9]), .ZN(n_24_33));
   NAND2_X1 i_24_43 (.A1(n_190), .A2(n_56), .ZN(n_24_34));
   NAND2_X1 i_24_44 (.A1(n_191), .A2(n_55), .ZN(n_24_35));
   NAND2_X1 i_24_45 (.A1(n_193), .A2(multiplicand[8]), .ZN(n_24_36));
   NAND4_X1 i_24_46 (.A1(n_24_33), .A2(n_24_34), .A3(n_24_35), .A4(n_24_36), 
      .ZN(n_203));
   NAND2_X1 i_24_47 (.A1(n_192), .A2(multiplicand[10]), .ZN(n_24_37));
   NAND2_X1 i_24_48 (.A1(n_190), .A2(n_57), .ZN(n_24_38));
   NAND2_X1 i_24_49 (.A1(n_191), .A2(n_56), .ZN(n_24_39));
   NAND2_X1 i_24_50 (.A1(n_193), .A2(multiplicand[9]), .ZN(n_24_40));
   NAND4_X1 i_24_51 (.A1(n_24_37), .A2(n_24_38), .A3(n_24_39), .A4(n_24_40), 
      .ZN(n_204));
   NAND2_X1 i_24_52 (.A1(n_192), .A2(multiplicand[11]), .ZN(n_24_41));
   NAND2_X1 i_24_53 (.A1(n_190), .A2(n_58), .ZN(n_24_42));
   NAND2_X1 i_24_54 (.A1(n_191), .A2(n_57), .ZN(n_24_43));
   NAND2_X1 i_24_55 (.A1(n_193), .A2(multiplicand[10]), .ZN(n_24_44));
   NAND4_X1 i_24_56 (.A1(n_24_41), .A2(n_24_42), .A3(n_24_43), .A4(n_24_44), 
      .ZN(n_205));
   NAND2_X1 i_24_57 (.A1(n_192), .A2(multiplicand[12]), .ZN(n_24_45));
   NAND2_X1 i_24_58 (.A1(n_190), .A2(n_59), .ZN(n_24_46));
   NAND2_X1 i_24_59 (.A1(n_191), .A2(n_58), .ZN(n_24_47));
   NAND2_X1 i_24_60 (.A1(n_193), .A2(multiplicand[11]), .ZN(n_24_48));
   NAND4_X1 i_24_61 (.A1(n_24_45), .A2(n_24_46), .A3(n_24_47), .A4(n_24_48), 
      .ZN(n_206));
   NAND2_X1 i_24_62 (.A1(n_192), .A2(multiplicand[13]), .ZN(n_24_49));
   NAND2_X1 i_24_63 (.A1(n_190), .A2(n_60), .ZN(n_24_50));
   NAND2_X1 i_24_64 (.A1(n_191), .A2(n_59), .ZN(n_24_51));
   NAND2_X1 i_24_65 (.A1(n_193), .A2(multiplicand[12]), .ZN(n_24_52));
   NAND4_X1 i_24_66 (.A1(n_24_49), .A2(n_24_50), .A3(n_24_51), .A4(n_24_52), 
      .ZN(n_207));
   NAND2_X1 i_24_67 (.A1(n_192), .A2(multiplicand[14]), .ZN(n_24_53));
   NAND2_X1 i_24_68 (.A1(n_190), .A2(n_61), .ZN(n_24_54));
   NAND2_X1 i_24_69 (.A1(n_191), .A2(n_60), .ZN(n_24_55));
   NAND2_X1 i_24_70 (.A1(n_193), .A2(multiplicand[13]), .ZN(n_24_56));
   NAND4_X1 i_24_71 (.A1(n_24_53), .A2(n_24_54), .A3(n_24_55), .A4(n_24_56), 
      .ZN(n_208));
   NAND2_X1 i_24_72 (.A1(n_192), .A2(multiplicand[15]), .ZN(n_24_57));
   NAND2_X1 i_24_73 (.A1(n_190), .A2(n_62), .ZN(n_24_58));
   NAND2_X1 i_24_74 (.A1(n_191), .A2(n_61), .ZN(n_24_59));
   NAND2_X1 i_24_75 (.A1(n_193), .A2(multiplicand[14]), .ZN(n_24_60));
   NAND4_X1 i_24_76 (.A1(n_24_57), .A2(n_24_58), .A3(n_24_59), .A4(n_24_60), 
      .ZN(n_209));
   NAND2_X1 i_24_77 (.A1(n_192), .A2(multiplicand[16]), .ZN(n_24_61));
   NAND2_X1 i_24_78 (.A1(n_190), .A2(n_63), .ZN(n_24_62));
   NAND2_X1 i_24_79 (.A1(n_191), .A2(n_62), .ZN(n_24_63));
   NAND2_X1 i_24_80 (.A1(n_193), .A2(multiplicand[15]), .ZN(n_24_64));
   NAND4_X1 i_24_81 (.A1(n_24_61), .A2(n_24_62), .A3(n_24_63), .A4(n_24_64), 
      .ZN(n_210));
   NAND2_X1 i_24_82 (.A1(n_192), .A2(multiplicand[17]), .ZN(n_24_65));
   NAND2_X1 i_24_83 (.A1(n_190), .A2(n_64), .ZN(n_24_66));
   NAND2_X1 i_24_84 (.A1(n_191), .A2(n_63), .ZN(n_24_67));
   NAND2_X1 i_24_85 (.A1(n_193), .A2(multiplicand[16]), .ZN(n_24_68));
   NAND4_X1 i_24_86 (.A1(n_24_65), .A2(n_24_66), .A3(n_24_67), .A4(n_24_68), 
      .ZN(n_211));
   NAND2_X1 i_24_87 (.A1(n_192), .A2(multiplicand[18]), .ZN(n_24_69));
   NAND2_X1 i_24_88 (.A1(n_190), .A2(n_65), .ZN(n_24_70));
   NAND2_X1 i_24_89 (.A1(n_191), .A2(n_64), .ZN(n_24_71));
   NAND2_X1 i_24_90 (.A1(n_193), .A2(multiplicand[17]), .ZN(n_24_72));
   NAND4_X1 i_24_91 (.A1(n_24_69), .A2(n_24_70), .A3(n_24_71), .A4(n_24_72), 
      .ZN(n_212));
   NAND2_X1 i_24_92 (.A1(n_192), .A2(multiplicand[19]), .ZN(n_24_73));
   NAND2_X1 i_24_93 (.A1(n_190), .A2(n_66), .ZN(n_24_74));
   NAND2_X1 i_24_94 (.A1(n_191), .A2(n_65), .ZN(n_24_75));
   NAND2_X1 i_24_95 (.A1(n_193), .A2(multiplicand[18]), .ZN(n_24_76));
   NAND4_X1 i_24_96 (.A1(n_24_73), .A2(n_24_74), .A3(n_24_75), .A4(n_24_76), 
      .ZN(n_213));
   NAND2_X1 i_24_97 (.A1(n_192), .A2(multiplicand[20]), .ZN(n_24_77));
   NAND2_X1 i_24_98 (.A1(n_190), .A2(n_67), .ZN(n_24_78));
   NAND2_X1 i_24_99 (.A1(n_191), .A2(n_66), .ZN(n_24_79));
   NAND2_X1 i_24_100 (.A1(n_193), .A2(multiplicand[19]), .ZN(n_24_80));
   NAND4_X1 i_24_101 (.A1(n_24_77), .A2(n_24_78), .A3(n_24_79), .A4(n_24_80), 
      .ZN(n_214));
   NAND2_X1 i_24_102 (.A1(n_192), .A2(multiplicand[21]), .ZN(n_24_81));
   NAND2_X1 i_24_103 (.A1(n_190), .A2(n_68), .ZN(n_24_82));
   NAND2_X1 i_24_104 (.A1(n_191), .A2(n_67), .ZN(n_24_83));
   NAND2_X1 i_24_105 (.A1(n_193), .A2(multiplicand[20]), .ZN(n_24_84));
   NAND4_X1 i_24_106 (.A1(n_24_81), .A2(n_24_82), .A3(n_24_83), .A4(n_24_84), 
      .ZN(n_215));
   NAND2_X1 i_24_107 (.A1(n_192), .A2(multiplicand[22]), .ZN(n_24_85));
   NAND2_X1 i_24_108 (.A1(n_190), .A2(n_69), .ZN(n_24_86));
   NAND2_X1 i_24_109 (.A1(n_191), .A2(n_68), .ZN(n_24_87));
   NAND2_X1 i_24_110 (.A1(n_193), .A2(multiplicand[21]), .ZN(n_24_88));
   NAND4_X1 i_24_111 (.A1(n_24_85), .A2(n_24_86), .A3(n_24_87), .A4(n_24_88), 
      .ZN(n_216));
   NAND2_X1 i_24_112 (.A1(n_192), .A2(multiplicand[23]), .ZN(n_24_89));
   NAND2_X1 i_24_113 (.A1(n_190), .A2(n_70), .ZN(n_24_90));
   NAND2_X1 i_24_114 (.A1(n_191), .A2(n_69), .ZN(n_24_91));
   NAND2_X1 i_24_115 (.A1(n_193), .A2(multiplicand[22]), .ZN(n_24_92));
   NAND4_X1 i_24_116 (.A1(n_24_89), .A2(n_24_90), .A3(n_24_91), .A4(n_24_92), 
      .ZN(n_217));
   NAND2_X1 i_24_117 (.A1(n_192), .A2(multiplicand[24]), .ZN(n_24_93));
   NAND2_X1 i_24_118 (.A1(n_190), .A2(n_71), .ZN(n_24_94));
   NAND2_X1 i_24_119 (.A1(n_191), .A2(n_70), .ZN(n_24_95));
   NAND2_X1 i_24_120 (.A1(n_193), .A2(multiplicand[23]), .ZN(n_24_96));
   NAND4_X1 i_24_121 (.A1(n_24_93), .A2(n_24_94), .A3(n_24_95), .A4(n_24_96), 
      .ZN(n_218));
   NAND2_X1 i_24_122 (.A1(n_192), .A2(multiplicand[25]), .ZN(n_24_97));
   NAND2_X1 i_24_123 (.A1(n_190), .A2(n_72), .ZN(n_24_98));
   NAND2_X1 i_24_124 (.A1(n_191), .A2(n_71), .ZN(n_24_99));
   NAND2_X1 i_24_125 (.A1(n_193), .A2(multiplicand[24]), .ZN(n_24_100));
   NAND4_X1 i_24_126 (.A1(n_24_97), .A2(n_24_98), .A3(n_24_99), .A4(n_24_100), 
      .ZN(n_219));
   NAND2_X1 i_24_127 (.A1(n_192), .A2(multiplicand[26]), .ZN(n_24_101));
   NAND2_X1 i_24_128 (.A1(n_190), .A2(n_73), .ZN(n_24_102));
   NAND2_X1 i_24_129 (.A1(n_191), .A2(n_72), .ZN(n_24_103));
   NAND2_X1 i_24_130 (.A1(n_193), .A2(multiplicand[25]), .ZN(n_24_104));
   NAND4_X1 i_24_131 (.A1(n_24_101), .A2(n_24_102), .A3(n_24_103), .A4(n_24_104), 
      .ZN(n_220));
   NAND2_X1 i_24_132 (.A1(n_192), .A2(multiplicand[27]), .ZN(n_24_105));
   NAND2_X1 i_24_133 (.A1(n_190), .A2(n_74), .ZN(n_24_106));
   NAND2_X1 i_24_134 (.A1(n_191), .A2(n_73), .ZN(n_24_107));
   NAND2_X1 i_24_135 (.A1(n_193), .A2(multiplicand[26]), .ZN(n_24_108));
   NAND4_X1 i_24_136 (.A1(n_24_105), .A2(n_24_106), .A3(n_24_107), .A4(n_24_108), 
      .ZN(n_221));
   NAND2_X1 i_24_137 (.A1(n_192), .A2(multiplicand[28]), .ZN(n_24_109));
   NAND2_X1 i_24_138 (.A1(n_190), .A2(n_75), .ZN(n_24_110));
   NAND2_X1 i_24_139 (.A1(n_191), .A2(n_74), .ZN(n_24_111));
   NAND2_X1 i_24_140 (.A1(n_193), .A2(multiplicand[27]), .ZN(n_24_112));
   NAND4_X1 i_24_141 (.A1(n_24_109), .A2(n_24_110), .A3(n_24_111), .A4(n_24_112), 
      .ZN(n_222));
   NAND2_X1 i_24_142 (.A1(n_192), .A2(multiplicand[29]), .ZN(n_24_113));
   NAND2_X1 i_24_143 (.A1(n_190), .A2(n_76), .ZN(n_24_114));
   NAND2_X1 i_24_144 (.A1(n_191), .A2(n_75), .ZN(n_24_115));
   NAND2_X1 i_24_145 (.A1(n_193), .A2(multiplicand[28]), .ZN(n_24_116));
   NAND4_X1 i_24_146 (.A1(n_24_113), .A2(n_24_114), .A3(n_24_115), .A4(n_24_116), 
      .ZN(n_223));
   NAND2_X1 i_24_147 (.A1(n_192), .A2(multiplicand[30]), .ZN(n_24_117));
   NAND2_X1 i_24_148 (.A1(n_190), .A2(n_77), .ZN(n_24_118));
   NAND2_X1 i_24_149 (.A1(n_191), .A2(n_76), .ZN(n_24_119));
   NAND2_X1 i_24_150 (.A1(n_193), .A2(multiplicand[29]), .ZN(n_24_120));
   NAND4_X1 i_24_151 (.A1(n_24_117), .A2(n_24_118), .A3(n_24_119), .A4(n_24_120), 
      .ZN(n_224));
   NAND2_X1 i_24_152 (.A1(n_192), .A2(multiplicand[31]), .ZN(n_24_121));
   NAND2_X1 i_24_153 (.A1(n_190), .A2(n_78), .ZN(n_24_122));
   NAND2_X1 i_24_154 (.A1(n_191), .A2(n_77), .ZN(n_24_123));
   NAND2_X1 i_24_155 (.A1(n_193), .A2(multiplicand[30]), .ZN(n_24_124));
   NAND4_X1 i_24_156 (.A1(n_24_121), .A2(n_24_122), .A3(n_24_123), .A4(n_24_124), 
      .ZN(n_225));
   NAND2_X1 i_24_157 (.A1(n_191), .A2(n_78), .ZN(n_24_125));
   NAND2_X1 i_24_158 (.A1(n_193), .A2(multiplicand[31]), .ZN(n_24_126));
   NAND4_X1 i_24_159 (.A1(n_24_121), .A2(n_24_122), .A3(n_24_125), .A4(n_24_126), 
      .ZN(n_226));
   INV_X1 i_25_0 (.A(n_12), .ZN(n_25_0));
   AND3_X1 i_25_1 (.A1(n_25_0), .A2(n_13), .A3(n_14), .ZN(n_227));
   INV_X1 i_25_2 (.A(n_13), .ZN(n_25_1));
   AND3_X1 i_25_3 (.A1(n_25_1), .A2(n_12), .A3(n_14), .ZN(n_228));
   NOR3_X1 i_25_4 (.A1(n_25_1), .A2(n_12), .A3(n_14), .ZN(n_229));
   NOR3_X1 i_25_5 (.A1(n_25_0), .A2(n_13), .A3(n_14), .ZN(n_230));
   AOI22_X1 i_26_0 (.A1(n_229), .A2(multiplicand[0]), .B1(n_227), .B2(
      multiplicand[0]), .ZN(n_26_0));
   INV_X1 i_26_1 (.A(n_26_0), .ZN(n_231));
   NAND2_X1 i_26_2 (.A1(n_229), .A2(multiplicand[1]), .ZN(n_26_1));
   NAND2_X1 i_26_3 (.A1(n_227), .A2(n_48), .ZN(n_26_2));
   NAND2_X1 i_26_4 (.A1(n_228), .A2(multiplicand[0]), .ZN(n_26_3));
   NAND2_X1 i_26_5 (.A1(n_230), .A2(multiplicand[0]), .ZN(n_26_4));
   NAND4_X1 i_26_6 (.A1(n_26_1), .A2(n_26_2), .A3(n_26_3), .A4(n_26_4), .ZN(
      n_232));
   NAND2_X1 i_26_7 (.A1(n_229), .A2(multiplicand[2]), .ZN(n_26_5));
   NAND2_X1 i_26_8 (.A1(n_227), .A2(n_49), .ZN(n_26_6));
   NAND2_X1 i_26_9 (.A1(n_228), .A2(n_48), .ZN(n_26_7));
   NAND2_X1 i_26_10 (.A1(n_230), .A2(multiplicand[1]), .ZN(n_26_8));
   NAND4_X1 i_26_11 (.A1(n_26_5), .A2(n_26_6), .A3(n_26_7), .A4(n_26_8), 
      .ZN(n_233));
   NAND2_X1 i_26_12 (.A1(n_229), .A2(multiplicand[3]), .ZN(n_26_9));
   NAND2_X1 i_26_13 (.A1(n_227), .A2(n_50), .ZN(n_26_10));
   NAND2_X1 i_26_14 (.A1(n_228), .A2(n_49), .ZN(n_26_11));
   NAND2_X1 i_26_15 (.A1(n_230), .A2(multiplicand[2]), .ZN(n_26_12));
   NAND4_X1 i_26_16 (.A1(n_26_9), .A2(n_26_10), .A3(n_26_11), .A4(n_26_12), 
      .ZN(n_234));
   NAND2_X1 i_26_17 (.A1(n_229), .A2(multiplicand[4]), .ZN(n_26_13));
   NAND2_X1 i_26_18 (.A1(n_227), .A2(n_51), .ZN(n_26_14));
   NAND2_X1 i_26_19 (.A1(n_228), .A2(n_50), .ZN(n_26_15));
   NAND2_X1 i_26_20 (.A1(n_230), .A2(multiplicand[3]), .ZN(n_26_16));
   NAND4_X1 i_26_21 (.A1(n_26_13), .A2(n_26_14), .A3(n_26_15), .A4(n_26_16), 
      .ZN(n_235));
   NAND2_X1 i_26_22 (.A1(n_229), .A2(multiplicand[5]), .ZN(n_26_17));
   NAND2_X1 i_26_23 (.A1(n_227), .A2(n_52), .ZN(n_26_18));
   NAND2_X1 i_26_24 (.A1(n_228), .A2(n_51), .ZN(n_26_19));
   NAND2_X1 i_26_25 (.A1(n_230), .A2(multiplicand[4]), .ZN(n_26_20));
   NAND4_X1 i_26_26 (.A1(n_26_17), .A2(n_26_18), .A3(n_26_19), .A4(n_26_20), 
      .ZN(n_236));
   NAND2_X1 i_26_27 (.A1(n_229), .A2(multiplicand[6]), .ZN(n_26_21));
   NAND2_X1 i_26_28 (.A1(n_227), .A2(n_53), .ZN(n_26_22));
   NAND2_X1 i_26_29 (.A1(n_228), .A2(n_52), .ZN(n_26_23));
   NAND2_X1 i_26_30 (.A1(n_230), .A2(multiplicand[5]), .ZN(n_26_24));
   NAND4_X1 i_26_31 (.A1(n_26_21), .A2(n_26_22), .A3(n_26_23), .A4(n_26_24), 
      .ZN(n_237));
   NAND2_X1 i_26_32 (.A1(n_229), .A2(multiplicand[7]), .ZN(n_26_25));
   NAND2_X1 i_26_33 (.A1(n_227), .A2(n_54), .ZN(n_26_26));
   NAND2_X1 i_26_34 (.A1(n_228), .A2(n_53), .ZN(n_26_27));
   NAND2_X1 i_26_35 (.A1(n_230), .A2(multiplicand[6]), .ZN(n_26_28));
   NAND4_X1 i_26_36 (.A1(n_26_25), .A2(n_26_26), .A3(n_26_27), .A4(n_26_28), 
      .ZN(n_238));
   NAND2_X1 i_26_37 (.A1(n_229), .A2(multiplicand[8]), .ZN(n_26_29));
   NAND2_X1 i_26_38 (.A1(n_227), .A2(n_55), .ZN(n_26_30));
   NAND2_X1 i_26_39 (.A1(n_228), .A2(n_54), .ZN(n_26_31));
   NAND2_X1 i_26_40 (.A1(n_230), .A2(multiplicand[7]), .ZN(n_26_32));
   NAND4_X1 i_26_41 (.A1(n_26_29), .A2(n_26_30), .A3(n_26_31), .A4(n_26_32), 
      .ZN(n_239));
   NAND2_X1 i_26_42 (.A1(n_229), .A2(multiplicand[9]), .ZN(n_26_33));
   NAND2_X1 i_26_43 (.A1(n_227), .A2(n_56), .ZN(n_26_34));
   NAND2_X1 i_26_44 (.A1(n_228), .A2(n_55), .ZN(n_26_35));
   NAND2_X1 i_26_45 (.A1(n_230), .A2(multiplicand[8]), .ZN(n_26_36));
   NAND4_X1 i_26_46 (.A1(n_26_33), .A2(n_26_34), .A3(n_26_35), .A4(n_26_36), 
      .ZN(n_240));
   NAND2_X1 i_26_47 (.A1(n_229), .A2(multiplicand[10]), .ZN(n_26_37));
   NAND2_X1 i_26_48 (.A1(n_227), .A2(n_57), .ZN(n_26_38));
   NAND2_X1 i_26_49 (.A1(n_228), .A2(n_56), .ZN(n_26_39));
   NAND2_X1 i_26_50 (.A1(n_230), .A2(multiplicand[9]), .ZN(n_26_40));
   NAND4_X1 i_26_51 (.A1(n_26_37), .A2(n_26_38), .A3(n_26_39), .A4(n_26_40), 
      .ZN(n_241));
   NAND2_X1 i_26_52 (.A1(n_229), .A2(multiplicand[11]), .ZN(n_26_41));
   NAND2_X1 i_26_53 (.A1(n_227), .A2(n_58), .ZN(n_26_42));
   NAND2_X1 i_26_54 (.A1(n_228), .A2(n_57), .ZN(n_26_43));
   NAND2_X1 i_26_55 (.A1(n_230), .A2(multiplicand[10]), .ZN(n_26_44));
   NAND4_X1 i_26_56 (.A1(n_26_41), .A2(n_26_42), .A3(n_26_43), .A4(n_26_44), 
      .ZN(n_242));
   NAND2_X1 i_26_57 (.A1(n_229), .A2(multiplicand[12]), .ZN(n_26_45));
   NAND2_X1 i_26_58 (.A1(n_227), .A2(n_59), .ZN(n_26_46));
   NAND2_X1 i_26_59 (.A1(n_228), .A2(n_58), .ZN(n_26_47));
   NAND2_X1 i_26_60 (.A1(n_230), .A2(multiplicand[11]), .ZN(n_26_48));
   NAND4_X1 i_26_61 (.A1(n_26_45), .A2(n_26_46), .A3(n_26_47), .A4(n_26_48), 
      .ZN(n_243));
   NAND2_X1 i_26_62 (.A1(n_229), .A2(multiplicand[13]), .ZN(n_26_49));
   NAND2_X1 i_26_63 (.A1(n_227), .A2(n_60), .ZN(n_26_50));
   NAND2_X1 i_26_64 (.A1(n_228), .A2(n_59), .ZN(n_26_51));
   NAND2_X1 i_26_65 (.A1(n_230), .A2(multiplicand[12]), .ZN(n_26_52));
   NAND4_X1 i_26_66 (.A1(n_26_49), .A2(n_26_50), .A3(n_26_51), .A4(n_26_52), 
      .ZN(n_244));
   NAND2_X1 i_26_67 (.A1(n_229), .A2(multiplicand[14]), .ZN(n_26_53));
   NAND2_X1 i_26_68 (.A1(n_227), .A2(n_61), .ZN(n_26_54));
   NAND2_X1 i_26_69 (.A1(n_228), .A2(n_60), .ZN(n_26_55));
   NAND2_X1 i_26_70 (.A1(n_230), .A2(multiplicand[13]), .ZN(n_26_56));
   NAND4_X1 i_26_71 (.A1(n_26_53), .A2(n_26_54), .A3(n_26_55), .A4(n_26_56), 
      .ZN(n_245));
   NAND2_X1 i_26_72 (.A1(n_229), .A2(multiplicand[15]), .ZN(n_26_57));
   NAND2_X1 i_26_73 (.A1(n_227), .A2(n_62), .ZN(n_26_58));
   NAND2_X1 i_26_74 (.A1(n_228), .A2(n_61), .ZN(n_26_59));
   NAND2_X1 i_26_75 (.A1(n_230), .A2(multiplicand[14]), .ZN(n_26_60));
   NAND4_X1 i_26_76 (.A1(n_26_57), .A2(n_26_58), .A3(n_26_59), .A4(n_26_60), 
      .ZN(n_246));
   NAND2_X1 i_26_77 (.A1(n_229), .A2(multiplicand[16]), .ZN(n_26_61));
   NAND2_X1 i_26_78 (.A1(n_227), .A2(n_63), .ZN(n_26_62));
   NAND2_X1 i_26_79 (.A1(n_228), .A2(n_62), .ZN(n_26_63));
   NAND2_X1 i_26_80 (.A1(n_230), .A2(multiplicand[15]), .ZN(n_26_64));
   NAND4_X1 i_26_81 (.A1(n_26_61), .A2(n_26_62), .A3(n_26_63), .A4(n_26_64), 
      .ZN(n_247));
   NAND2_X1 i_26_82 (.A1(n_229), .A2(multiplicand[17]), .ZN(n_26_65));
   NAND2_X1 i_26_83 (.A1(n_227), .A2(n_64), .ZN(n_26_66));
   NAND2_X1 i_26_84 (.A1(n_228), .A2(n_63), .ZN(n_26_67));
   NAND2_X1 i_26_85 (.A1(n_230), .A2(multiplicand[16]), .ZN(n_26_68));
   NAND4_X1 i_26_86 (.A1(n_26_65), .A2(n_26_66), .A3(n_26_67), .A4(n_26_68), 
      .ZN(n_248));
   NAND2_X1 i_26_87 (.A1(n_229), .A2(multiplicand[18]), .ZN(n_26_69));
   NAND2_X1 i_26_88 (.A1(n_227), .A2(n_65), .ZN(n_26_70));
   NAND2_X1 i_26_89 (.A1(n_228), .A2(n_64), .ZN(n_26_71));
   NAND2_X1 i_26_90 (.A1(n_230), .A2(multiplicand[17]), .ZN(n_26_72));
   NAND4_X1 i_26_91 (.A1(n_26_69), .A2(n_26_70), .A3(n_26_71), .A4(n_26_72), 
      .ZN(n_249));
   NAND2_X1 i_26_92 (.A1(n_229), .A2(multiplicand[19]), .ZN(n_26_73));
   NAND2_X1 i_26_93 (.A1(n_227), .A2(n_66), .ZN(n_26_74));
   NAND2_X1 i_26_94 (.A1(n_228), .A2(n_65), .ZN(n_26_75));
   NAND2_X1 i_26_95 (.A1(n_230), .A2(multiplicand[18]), .ZN(n_26_76));
   NAND4_X1 i_26_96 (.A1(n_26_73), .A2(n_26_74), .A3(n_26_75), .A4(n_26_76), 
      .ZN(n_250));
   NAND2_X1 i_26_97 (.A1(n_229), .A2(multiplicand[20]), .ZN(n_26_77));
   NAND2_X1 i_26_98 (.A1(n_227), .A2(n_67), .ZN(n_26_78));
   NAND2_X1 i_26_99 (.A1(n_228), .A2(n_66), .ZN(n_26_79));
   NAND2_X1 i_26_100 (.A1(n_230), .A2(multiplicand[19]), .ZN(n_26_80));
   NAND4_X1 i_26_101 (.A1(n_26_77), .A2(n_26_78), .A3(n_26_79), .A4(n_26_80), 
      .ZN(n_251));
   NAND2_X1 i_26_102 (.A1(n_229), .A2(multiplicand[21]), .ZN(n_26_81));
   NAND2_X1 i_26_103 (.A1(n_227), .A2(n_68), .ZN(n_26_82));
   NAND2_X1 i_26_104 (.A1(n_228), .A2(n_67), .ZN(n_26_83));
   NAND2_X1 i_26_105 (.A1(n_230), .A2(multiplicand[20]), .ZN(n_26_84));
   NAND4_X1 i_26_106 (.A1(n_26_81), .A2(n_26_82), .A3(n_26_83), .A4(n_26_84), 
      .ZN(n_252));
   NAND2_X1 i_26_107 (.A1(n_229), .A2(multiplicand[22]), .ZN(n_26_85));
   NAND2_X1 i_26_108 (.A1(n_227), .A2(n_69), .ZN(n_26_86));
   NAND2_X1 i_26_109 (.A1(n_228), .A2(n_68), .ZN(n_26_87));
   NAND2_X1 i_26_110 (.A1(n_230), .A2(multiplicand[21]), .ZN(n_26_88));
   NAND4_X1 i_26_111 (.A1(n_26_85), .A2(n_26_86), .A3(n_26_87), .A4(n_26_88), 
      .ZN(n_253));
   NAND2_X1 i_26_112 (.A1(n_229), .A2(multiplicand[23]), .ZN(n_26_89));
   NAND2_X1 i_26_113 (.A1(n_227), .A2(n_70), .ZN(n_26_90));
   NAND2_X1 i_26_114 (.A1(n_228), .A2(n_69), .ZN(n_26_91));
   NAND2_X1 i_26_115 (.A1(n_230), .A2(multiplicand[22]), .ZN(n_26_92));
   NAND4_X1 i_26_116 (.A1(n_26_89), .A2(n_26_90), .A3(n_26_91), .A4(n_26_92), 
      .ZN(n_254));
   NAND2_X1 i_26_117 (.A1(n_229), .A2(multiplicand[24]), .ZN(n_26_93));
   NAND2_X1 i_26_118 (.A1(n_227), .A2(n_71), .ZN(n_26_94));
   NAND2_X1 i_26_119 (.A1(n_228), .A2(n_70), .ZN(n_26_95));
   NAND2_X1 i_26_120 (.A1(n_230), .A2(multiplicand[23]), .ZN(n_26_96));
   NAND4_X1 i_26_121 (.A1(n_26_93), .A2(n_26_94), .A3(n_26_95), .A4(n_26_96), 
      .ZN(n_255));
   NAND2_X1 i_26_122 (.A1(n_229), .A2(multiplicand[25]), .ZN(n_26_97));
   NAND2_X1 i_26_123 (.A1(n_227), .A2(n_72), .ZN(n_26_98));
   NAND2_X1 i_26_124 (.A1(n_228), .A2(n_71), .ZN(n_26_99));
   NAND2_X1 i_26_125 (.A1(n_230), .A2(multiplicand[24]), .ZN(n_26_100));
   NAND4_X1 i_26_126 (.A1(n_26_97), .A2(n_26_98), .A3(n_26_99), .A4(n_26_100), 
      .ZN(n_256));
   NAND2_X1 i_26_127 (.A1(n_229), .A2(multiplicand[26]), .ZN(n_26_101));
   NAND2_X1 i_26_128 (.A1(n_227), .A2(n_73), .ZN(n_26_102));
   NAND2_X1 i_26_129 (.A1(n_228), .A2(n_72), .ZN(n_26_103));
   NAND2_X1 i_26_130 (.A1(n_230), .A2(multiplicand[25]), .ZN(n_26_104));
   NAND4_X1 i_26_131 (.A1(n_26_101), .A2(n_26_102), .A3(n_26_103), .A4(n_26_104), 
      .ZN(n_257));
   NAND2_X1 i_26_132 (.A1(n_229), .A2(multiplicand[27]), .ZN(n_26_105));
   NAND2_X1 i_26_133 (.A1(n_227), .A2(n_74), .ZN(n_26_106));
   NAND2_X1 i_26_134 (.A1(n_228), .A2(n_73), .ZN(n_26_107));
   NAND2_X1 i_26_135 (.A1(n_230), .A2(multiplicand[26]), .ZN(n_26_108));
   NAND4_X1 i_26_136 (.A1(n_26_105), .A2(n_26_106), .A3(n_26_107), .A4(n_26_108), 
      .ZN(n_258));
   NAND2_X1 i_26_137 (.A1(n_229), .A2(multiplicand[28]), .ZN(n_26_109));
   NAND2_X1 i_26_138 (.A1(n_227), .A2(n_75), .ZN(n_26_110));
   NAND2_X1 i_26_139 (.A1(n_228), .A2(n_74), .ZN(n_26_111));
   NAND2_X1 i_26_140 (.A1(n_230), .A2(multiplicand[27]), .ZN(n_26_112));
   NAND4_X1 i_26_141 (.A1(n_26_109), .A2(n_26_110), .A3(n_26_111), .A4(n_26_112), 
      .ZN(n_259));
   NAND2_X1 i_26_142 (.A1(n_229), .A2(multiplicand[29]), .ZN(n_26_113));
   NAND2_X1 i_26_143 (.A1(n_227), .A2(n_76), .ZN(n_26_114));
   NAND2_X1 i_26_144 (.A1(n_228), .A2(n_75), .ZN(n_26_115));
   NAND2_X1 i_26_145 (.A1(n_230), .A2(multiplicand[28]), .ZN(n_26_116));
   NAND4_X1 i_26_146 (.A1(n_26_113), .A2(n_26_114), .A3(n_26_115), .A4(n_26_116), 
      .ZN(n_260));
   NAND2_X1 i_26_147 (.A1(n_229), .A2(multiplicand[30]), .ZN(n_26_117));
   NAND2_X1 i_26_148 (.A1(n_227), .A2(n_77), .ZN(n_26_118));
   NAND2_X1 i_26_149 (.A1(n_228), .A2(n_76), .ZN(n_26_119));
   NAND2_X1 i_26_150 (.A1(n_230), .A2(multiplicand[29]), .ZN(n_26_120));
   NAND4_X1 i_26_151 (.A1(n_26_117), .A2(n_26_118), .A3(n_26_119), .A4(n_26_120), 
      .ZN(n_261));
   NAND2_X1 i_26_152 (.A1(n_229), .A2(multiplicand[31]), .ZN(n_26_121));
   NAND2_X1 i_26_153 (.A1(n_227), .A2(n_78), .ZN(n_26_122));
   NAND2_X1 i_26_154 (.A1(n_228), .A2(n_77), .ZN(n_26_123));
   NAND2_X1 i_26_155 (.A1(n_230), .A2(multiplicand[30]), .ZN(n_26_124));
   NAND4_X1 i_26_156 (.A1(n_26_121), .A2(n_26_122), .A3(n_26_123), .A4(n_26_124), 
      .ZN(n_262));
   NAND2_X1 i_26_157 (.A1(n_228), .A2(n_78), .ZN(n_26_125));
   NAND2_X1 i_26_158 (.A1(n_230), .A2(multiplicand[31]), .ZN(n_26_126));
   NAND4_X1 i_26_159 (.A1(n_26_121), .A2(n_26_122), .A3(n_26_125), .A4(n_26_126), 
      .ZN(n_263));
   INV_X1 i_27_0 (.A(n_15), .ZN(n_27_0));
   AND3_X1 i_27_1 (.A1(n_27_0), .A2(n_16), .A3(n_17), .ZN(n_264));
   INV_X1 i_27_2 (.A(n_16), .ZN(n_27_1));
   AND3_X1 i_27_3 (.A1(n_27_1), .A2(n_15), .A3(n_17), .ZN(n_265));
   NOR3_X1 i_27_4 (.A1(n_27_1), .A2(n_15), .A3(n_17), .ZN(n_266));
   NOR3_X1 i_27_5 (.A1(n_27_0), .A2(n_16), .A3(n_17), .ZN(n_267));
   AOI22_X1 i_28_0 (.A1(n_266), .A2(multiplicand[0]), .B1(n_264), .B2(
      multiplicand[0]), .ZN(n_28_0));
   INV_X1 i_28_1 (.A(n_28_0), .ZN(n_268));
   NAND2_X1 i_28_2 (.A1(n_266), .A2(multiplicand[1]), .ZN(n_28_1));
   NAND2_X1 i_28_3 (.A1(n_264), .A2(n_48), .ZN(n_28_2));
   NAND2_X1 i_28_4 (.A1(n_265), .A2(multiplicand[0]), .ZN(n_28_3));
   NAND2_X1 i_28_5 (.A1(n_267), .A2(multiplicand[0]), .ZN(n_28_4));
   NAND4_X1 i_28_6 (.A1(n_28_1), .A2(n_28_2), .A3(n_28_3), .A4(n_28_4), .ZN(
      n_269));
   NAND2_X1 i_28_7 (.A1(n_266), .A2(multiplicand[2]), .ZN(n_28_5));
   NAND2_X1 i_28_8 (.A1(n_264), .A2(n_49), .ZN(n_28_6));
   NAND2_X1 i_28_9 (.A1(n_265), .A2(n_48), .ZN(n_28_7));
   NAND2_X1 i_28_10 (.A1(n_267), .A2(multiplicand[1]), .ZN(n_28_8));
   NAND4_X1 i_28_11 (.A1(n_28_5), .A2(n_28_6), .A3(n_28_7), .A4(n_28_8), 
      .ZN(n_270));
   NAND2_X1 i_28_12 (.A1(n_266), .A2(multiplicand[3]), .ZN(n_28_9));
   NAND2_X1 i_28_13 (.A1(n_264), .A2(n_50), .ZN(n_28_10));
   NAND2_X1 i_28_14 (.A1(n_265), .A2(n_49), .ZN(n_28_11));
   NAND2_X1 i_28_15 (.A1(n_267), .A2(multiplicand[2]), .ZN(n_28_12));
   NAND4_X1 i_28_16 (.A1(n_28_9), .A2(n_28_10), .A3(n_28_11), .A4(n_28_12), 
      .ZN(n_271));
   NAND2_X1 i_28_17 (.A1(n_266), .A2(multiplicand[4]), .ZN(n_28_13));
   NAND2_X1 i_28_18 (.A1(n_264), .A2(n_51), .ZN(n_28_14));
   NAND2_X1 i_28_19 (.A1(n_265), .A2(n_50), .ZN(n_28_15));
   NAND2_X1 i_28_20 (.A1(n_267), .A2(multiplicand[3]), .ZN(n_28_16));
   NAND4_X1 i_28_21 (.A1(n_28_13), .A2(n_28_14), .A3(n_28_15), .A4(n_28_16), 
      .ZN(n_272));
   NAND2_X1 i_28_22 (.A1(n_266), .A2(multiplicand[5]), .ZN(n_28_17));
   NAND2_X1 i_28_23 (.A1(n_264), .A2(n_52), .ZN(n_28_18));
   NAND2_X1 i_28_24 (.A1(n_265), .A2(n_51), .ZN(n_28_19));
   NAND2_X1 i_28_25 (.A1(n_267), .A2(multiplicand[4]), .ZN(n_28_20));
   NAND4_X1 i_28_26 (.A1(n_28_17), .A2(n_28_18), .A3(n_28_19), .A4(n_28_20), 
      .ZN(n_273));
   NAND2_X1 i_28_27 (.A1(n_266), .A2(multiplicand[6]), .ZN(n_28_21));
   NAND2_X1 i_28_28 (.A1(n_264), .A2(n_53), .ZN(n_28_22));
   NAND2_X1 i_28_29 (.A1(n_265), .A2(n_52), .ZN(n_28_23));
   NAND2_X1 i_28_30 (.A1(n_267), .A2(multiplicand[5]), .ZN(n_28_24));
   NAND4_X1 i_28_31 (.A1(n_28_21), .A2(n_28_22), .A3(n_28_23), .A4(n_28_24), 
      .ZN(n_274));
   NAND2_X1 i_28_32 (.A1(n_266), .A2(multiplicand[7]), .ZN(n_28_25));
   NAND2_X1 i_28_33 (.A1(n_264), .A2(n_54), .ZN(n_28_26));
   NAND2_X1 i_28_34 (.A1(n_265), .A2(n_53), .ZN(n_28_27));
   NAND2_X1 i_28_35 (.A1(n_267), .A2(multiplicand[6]), .ZN(n_28_28));
   NAND4_X1 i_28_36 (.A1(n_28_25), .A2(n_28_26), .A3(n_28_27), .A4(n_28_28), 
      .ZN(n_275));
   NAND2_X1 i_28_37 (.A1(n_266), .A2(multiplicand[8]), .ZN(n_28_29));
   NAND2_X1 i_28_38 (.A1(n_264), .A2(n_55), .ZN(n_28_30));
   NAND2_X1 i_28_39 (.A1(n_265), .A2(n_54), .ZN(n_28_31));
   NAND2_X1 i_28_40 (.A1(n_267), .A2(multiplicand[7]), .ZN(n_28_32));
   NAND4_X1 i_28_41 (.A1(n_28_29), .A2(n_28_30), .A3(n_28_31), .A4(n_28_32), 
      .ZN(n_276));
   NAND2_X1 i_28_42 (.A1(n_266), .A2(multiplicand[9]), .ZN(n_28_33));
   NAND2_X1 i_28_43 (.A1(n_264), .A2(n_56), .ZN(n_28_34));
   NAND2_X1 i_28_44 (.A1(n_265), .A2(n_55), .ZN(n_28_35));
   NAND2_X1 i_28_45 (.A1(n_267), .A2(multiplicand[8]), .ZN(n_28_36));
   NAND4_X1 i_28_46 (.A1(n_28_33), .A2(n_28_34), .A3(n_28_35), .A4(n_28_36), 
      .ZN(n_277));
   NAND2_X1 i_28_47 (.A1(n_266), .A2(multiplicand[10]), .ZN(n_28_37));
   NAND2_X1 i_28_48 (.A1(n_264), .A2(n_57), .ZN(n_28_38));
   NAND2_X1 i_28_49 (.A1(n_265), .A2(n_56), .ZN(n_28_39));
   NAND2_X1 i_28_50 (.A1(n_267), .A2(multiplicand[9]), .ZN(n_28_40));
   NAND4_X1 i_28_51 (.A1(n_28_37), .A2(n_28_38), .A3(n_28_39), .A4(n_28_40), 
      .ZN(n_278));
   NAND2_X1 i_28_52 (.A1(n_266), .A2(multiplicand[11]), .ZN(n_28_41));
   NAND2_X1 i_28_53 (.A1(n_264), .A2(n_58), .ZN(n_28_42));
   NAND2_X1 i_28_54 (.A1(n_265), .A2(n_57), .ZN(n_28_43));
   NAND2_X1 i_28_55 (.A1(n_267), .A2(multiplicand[10]), .ZN(n_28_44));
   NAND4_X1 i_28_56 (.A1(n_28_41), .A2(n_28_42), .A3(n_28_43), .A4(n_28_44), 
      .ZN(n_279));
   NAND2_X1 i_28_57 (.A1(n_266), .A2(multiplicand[12]), .ZN(n_28_45));
   NAND2_X1 i_28_58 (.A1(n_264), .A2(n_59), .ZN(n_28_46));
   NAND2_X1 i_28_59 (.A1(n_265), .A2(n_58), .ZN(n_28_47));
   NAND2_X1 i_28_60 (.A1(n_267), .A2(multiplicand[11]), .ZN(n_28_48));
   NAND4_X1 i_28_61 (.A1(n_28_45), .A2(n_28_46), .A3(n_28_47), .A4(n_28_48), 
      .ZN(n_280));
   NAND2_X1 i_28_62 (.A1(n_266), .A2(multiplicand[13]), .ZN(n_28_49));
   NAND2_X1 i_28_63 (.A1(n_264), .A2(n_60), .ZN(n_28_50));
   NAND2_X1 i_28_64 (.A1(n_265), .A2(n_59), .ZN(n_28_51));
   NAND2_X1 i_28_65 (.A1(n_267), .A2(multiplicand[12]), .ZN(n_28_52));
   NAND4_X1 i_28_66 (.A1(n_28_49), .A2(n_28_50), .A3(n_28_51), .A4(n_28_52), 
      .ZN(n_281));
   NAND2_X1 i_28_67 (.A1(n_266), .A2(multiplicand[14]), .ZN(n_28_53));
   NAND2_X1 i_28_68 (.A1(n_264), .A2(n_61), .ZN(n_28_54));
   NAND2_X1 i_28_69 (.A1(n_265), .A2(n_60), .ZN(n_28_55));
   NAND2_X1 i_28_70 (.A1(n_267), .A2(multiplicand[13]), .ZN(n_28_56));
   NAND4_X1 i_28_71 (.A1(n_28_53), .A2(n_28_54), .A3(n_28_55), .A4(n_28_56), 
      .ZN(n_282));
   NAND2_X1 i_28_72 (.A1(n_266), .A2(multiplicand[15]), .ZN(n_28_57));
   NAND2_X1 i_28_73 (.A1(n_264), .A2(n_62), .ZN(n_28_58));
   NAND2_X1 i_28_74 (.A1(n_265), .A2(n_61), .ZN(n_28_59));
   NAND2_X1 i_28_75 (.A1(n_267), .A2(multiplicand[14]), .ZN(n_28_60));
   NAND4_X1 i_28_76 (.A1(n_28_57), .A2(n_28_58), .A3(n_28_59), .A4(n_28_60), 
      .ZN(n_283));
   NAND2_X1 i_28_77 (.A1(n_266), .A2(multiplicand[16]), .ZN(n_28_61));
   NAND2_X1 i_28_78 (.A1(n_264), .A2(n_63), .ZN(n_28_62));
   NAND2_X1 i_28_79 (.A1(n_265), .A2(n_62), .ZN(n_28_63));
   NAND2_X1 i_28_80 (.A1(n_267), .A2(multiplicand[15]), .ZN(n_28_64));
   NAND4_X1 i_28_81 (.A1(n_28_61), .A2(n_28_62), .A3(n_28_63), .A4(n_28_64), 
      .ZN(n_284));
   NAND2_X1 i_28_82 (.A1(n_266), .A2(multiplicand[17]), .ZN(n_28_65));
   NAND2_X1 i_28_83 (.A1(n_264), .A2(n_64), .ZN(n_28_66));
   NAND2_X1 i_28_84 (.A1(n_265), .A2(n_63), .ZN(n_28_67));
   NAND2_X1 i_28_85 (.A1(n_267), .A2(multiplicand[16]), .ZN(n_28_68));
   NAND4_X1 i_28_86 (.A1(n_28_65), .A2(n_28_66), .A3(n_28_67), .A4(n_28_68), 
      .ZN(n_285));
   NAND2_X1 i_28_87 (.A1(n_266), .A2(multiplicand[18]), .ZN(n_28_69));
   NAND2_X1 i_28_88 (.A1(n_264), .A2(n_65), .ZN(n_28_70));
   NAND2_X1 i_28_89 (.A1(n_265), .A2(n_64), .ZN(n_28_71));
   NAND2_X1 i_28_90 (.A1(n_267), .A2(multiplicand[17]), .ZN(n_28_72));
   NAND4_X1 i_28_91 (.A1(n_28_69), .A2(n_28_70), .A3(n_28_71), .A4(n_28_72), 
      .ZN(n_286));
   NAND2_X1 i_28_92 (.A1(n_266), .A2(multiplicand[19]), .ZN(n_28_73));
   NAND2_X1 i_28_93 (.A1(n_264), .A2(n_66), .ZN(n_28_74));
   NAND2_X1 i_28_94 (.A1(n_265), .A2(n_65), .ZN(n_28_75));
   NAND2_X1 i_28_95 (.A1(n_267), .A2(multiplicand[18]), .ZN(n_28_76));
   NAND4_X1 i_28_96 (.A1(n_28_73), .A2(n_28_74), .A3(n_28_75), .A4(n_28_76), 
      .ZN(n_287));
   NAND2_X1 i_28_97 (.A1(n_266), .A2(multiplicand[20]), .ZN(n_28_77));
   NAND2_X1 i_28_98 (.A1(n_264), .A2(n_67), .ZN(n_28_78));
   NAND2_X1 i_28_99 (.A1(n_265), .A2(n_66), .ZN(n_28_79));
   NAND2_X1 i_28_100 (.A1(n_267), .A2(multiplicand[19]), .ZN(n_28_80));
   NAND4_X1 i_28_101 (.A1(n_28_77), .A2(n_28_78), .A3(n_28_79), .A4(n_28_80), 
      .ZN(n_288));
   NAND2_X1 i_28_102 (.A1(n_266), .A2(multiplicand[21]), .ZN(n_28_81));
   NAND2_X1 i_28_103 (.A1(n_264), .A2(n_68), .ZN(n_28_82));
   NAND2_X1 i_28_104 (.A1(n_265), .A2(n_67), .ZN(n_28_83));
   NAND2_X1 i_28_105 (.A1(n_267), .A2(multiplicand[20]), .ZN(n_28_84));
   NAND4_X1 i_28_106 (.A1(n_28_81), .A2(n_28_82), .A3(n_28_83), .A4(n_28_84), 
      .ZN(n_289));
   NAND2_X1 i_28_107 (.A1(n_266), .A2(multiplicand[22]), .ZN(n_28_85));
   NAND2_X1 i_28_108 (.A1(n_264), .A2(n_69), .ZN(n_28_86));
   NAND2_X1 i_28_109 (.A1(n_265), .A2(n_68), .ZN(n_28_87));
   NAND2_X1 i_28_110 (.A1(n_267), .A2(multiplicand[21]), .ZN(n_28_88));
   NAND4_X1 i_28_111 (.A1(n_28_85), .A2(n_28_86), .A3(n_28_87), .A4(n_28_88), 
      .ZN(n_290));
   NAND2_X1 i_28_112 (.A1(n_266), .A2(multiplicand[23]), .ZN(n_28_89));
   NAND2_X1 i_28_113 (.A1(n_264), .A2(n_70), .ZN(n_28_90));
   NAND2_X1 i_28_114 (.A1(n_265), .A2(n_69), .ZN(n_28_91));
   NAND2_X1 i_28_115 (.A1(n_267), .A2(multiplicand[22]), .ZN(n_28_92));
   NAND4_X1 i_28_116 (.A1(n_28_89), .A2(n_28_90), .A3(n_28_91), .A4(n_28_92), 
      .ZN(n_291));
   NAND2_X1 i_28_117 (.A1(n_266), .A2(multiplicand[24]), .ZN(n_28_93));
   NAND2_X1 i_28_118 (.A1(n_264), .A2(n_71), .ZN(n_28_94));
   NAND2_X1 i_28_119 (.A1(n_265), .A2(n_70), .ZN(n_28_95));
   NAND2_X1 i_28_120 (.A1(n_267), .A2(multiplicand[23]), .ZN(n_28_96));
   NAND4_X1 i_28_121 (.A1(n_28_93), .A2(n_28_94), .A3(n_28_95), .A4(n_28_96), 
      .ZN(n_292));
   NAND2_X1 i_28_122 (.A1(n_266), .A2(multiplicand[25]), .ZN(n_28_97));
   NAND2_X1 i_28_123 (.A1(n_264), .A2(n_72), .ZN(n_28_98));
   NAND2_X1 i_28_124 (.A1(n_265), .A2(n_71), .ZN(n_28_99));
   NAND2_X1 i_28_125 (.A1(n_267), .A2(multiplicand[24]), .ZN(n_28_100));
   NAND4_X1 i_28_126 (.A1(n_28_97), .A2(n_28_98), .A3(n_28_99), .A4(n_28_100), 
      .ZN(n_293));
   NAND2_X1 i_28_127 (.A1(n_266), .A2(multiplicand[26]), .ZN(n_28_101));
   NAND2_X1 i_28_128 (.A1(n_264), .A2(n_73), .ZN(n_28_102));
   NAND2_X1 i_28_129 (.A1(n_265), .A2(n_72), .ZN(n_28_103));
   NAND2_X1 i_28_130 (.A1(n_267), .A2(multiplicand[25]), .ZN(n_28_104));
   NAND4_X1 i_28_131 (.A1(n_28_101), .A2(n_28_102), .A3(n_28_103), .A4(n_28_104), 
      .ZN(n_294));
   NAND2_X1 i_28_132 (.A1(n_266), .A2(multiplicand[27]), .ZN(n_28_105));
   NAND2_X1 i_28_133 (.A1(n_264), .A2(n_74), .ZN(n_28_106));
   NAND2_X1 i_28_134 (.A1(n_265), .A2(n_73), .ZN(n_28_107));
   NAND2_X1 i_28_135 (.A1(n_267), .A2(multiplicand[26]), .ZN(n_28_108));
   NAND4_X1 i_28_136 (.A1(n_28_105), .A2(n_28_106), .A3(n_28_107), .A4(n_28_108), 
      .ZN(n_295));
   NAND2_X1 i_28_137 (.A1(n_266), .A2(multiplicand[28]), .ZN(n_28_109));
   NAND2_X1 i_28_138 (.A1(n_264), .A2(n_75), .ZN(n_28_110));
   NAND2_X1 i_28_139 (.A1(n_265), .A2(n_74), .ZN(n_28_111));
   NAND2_X1 i_28_140 (.A1(n_267), .A2(multiplicand[27]), .ZN(n_28_112));
   NAND4_X1 i_28_141 (.A1(n_28_109), .A2(n_28_110), .A3(n_28_111), .A4(n_28_112), 
      .ZN(n_296));
   NAND2_X1 i_28_142 (.A1(n_266), .A2(multiplicand[29]), .ZN(n_28_113));
   NAND2_X1 i_28_143 (.A1(n_264), .A2(n_76), .ZN(n_28_114));
   NAND2_X1 i_28_144 (.A1(n_265), .A2(n_75), .ZN(n_28_115));
   NAND2_X1 i_28_145 (.A1(n_267), .A2(multiplicand[28]), .ZN(n_28_116));
   NAND4_X1 i_28_146 (.A1(n_28_113), .A2(n_28_114), .A3(n_28_115), .A4(n_28_116), 
      .ZN(n_297));
   NAND2_X1 i_28_147 (.A1(n_266), .A2(multiplicand[30]), .ZN(n_28_117));
   NAND2_X1 i_28_148 (.A1(n_264), .A2(n_77), .ZN(n_28_118));
   NAND2_X1 i_28_149 (.A1(n_265), .A2(n_76), .ZN(n_28_119));
   NAND2_X1 i_28_150 (.A1(n_267), .A2(multiplicand[29]), .ZN(n_28_120));
   NAND4_X1 i_28_151 (.A1(n_28_117), .A2(n_28_118), .A3(n_28_119), .A4(n_28_120), 
      .ZN(n_298));
   NAND2_X1 i_28_152 (.A1(n_266), .A2(multiplicand[31]), .ZN(n_28_121));
   NAND2_X1 i_28_153 (.A1(n_264), .A2(n_78), .ZN(n_28_122));
   NAND2_X1 i_28_154 (.A1(n_265), .A2(n_77), .ZN(n_28_123));
   NAND2_X1 i_28_155 (.A1(n_267), .A2(multiplicand[30]), .ZN(n_28_124));
   NAND4_X1 i_28_156 (.A1(n_28_121), .A2(n_28_122), .A3(n_28_123), .A4(n_28_124), 
      .ZN(n_299));
   NAND2_X1 i_28_157 (.A1(n_265), .A2(n_78), .ZN(n_28_125));
   NAND2_X1 i_28_158 (.A1(n_267), .A2(multiplicand[31]), .ZN(n_28_126));
   NAND4_X1 i_28_159 (.A1(n_28_121), .A2(n_28_122), .A3(n_28_125), .A4(n_28_126), 
      .ZN(n_300));
   INV_X1 i_29_0 (.A(n_18), .ZN(n_29_0));
   AND3_X1 i_29_1 (.A1(n_29_0), .A2(n_19), .A3(n_20), .ZN(n_301));
   INV_X1 i_29_2 (.A(n_19), .ZN(n_29_1));
   AND3_X1 i_29_3 (.A1(n_29_1), .A2(n_18), .A3(n_20), .ZN(n_302));
   NOR3_X1 i_29_4 (.A1(n_29_1), .A2(n_18), .A3(n_20), .ZN(n_303));
   NOR3_X1 i_29_5 (.A1(n_29_0), .A2(n_19), .A3(n_20), .ZN(n_304));
   AOI22_X1 i_30_0 (.A1(n_303), .A2(multiplicand[0]), .B1(n_301), .B2(
      multiplicand[0]), .ZN(n_30_0));
   INV_X1 i_30_1 (.A(n_30_0), .ZN(n_305));
   NAND2_X1 i_30_2 (.A1(n_303), .A2(multiplicand[1]), .ZN(n_30_1));
   NAND2_X1 i_30_3 (.A1(n_301), .A2(n_48), .ZN(n_30_2));
   NAND2_X1 i_30_4 (.A1(n_302), .A2(multiplicand[0]), .ZN(n_30_3));
   NAND2_X1 i_30_5 (.A1(n_304), .A2(multiplicand[0]), .ZN(n_30_4));
   NAND4_X1 i_30_6 (.A1(n_30_1), .A2(n_30_2), .A3(n_30_3), .A4(n_30_4), .ZN(
      n_306));
   NAND2_X1 i_30_7 (.A1(n_303), .A2(multiplicand[2]), .ZN(n_30_5));
   NAND2_X1 i_30_8 (.A1(n_301), .A2(n_49), .ZN(n_30_6));
   NAND2_X1 i_30_9 (.A1(n_302), .A2(n_48), .ZN(n_30_7));
   NAND2_X1 i_30_10 (.A1(n_304), .A2(multiplicand[1]), .ZN(n_30_8));
   NAND4_X1 i_30_11 (.A1(n_30_5), .A2(n_30_6), .A3(n_30_7), .A4(n_30_8), 
      .ZN(n_307));
   NAND2_X1 i_30_12 (.A1(n_303), .A2(multiplicand[3]), .ZN(n_30_9));
   NAND2_X1 i_30_13 (.A1(n_301), .A2(n_50), .ZN(n_30_10));
   NAND2_X1 i_30_14 (.A1(n_302), .A2(n_49), .ZN(n_30_11));
   NAND2_X1 i_30_15 (.A1(n_304), .A2(multiplicand[2]), .ZN(n_30_12));
   NAND4_X1 i_30_16 (.A1(n_30_9), .A2(n_30_10), .A3(n_30_11), .A4(n_30_12), 
      .ZN(n_308));
   NAND2_X1 i_30_17 (.A1(n_303), .A2(multiplicand[4]), .ZN(n_30_13));
   NAND2_X1 i_30_18 (.A1(n_301), .A2(n_51), .ZN(n_30_14));
   NAND2_X1 i_30_19 (.A1(n_302), .A2(n_50), .ZN(n_30_15));
   NAND2_X1 i_30_20 (.A1(n_304), .A2(multiplicand[3]), .ZN(n_30_16));
   NAND4_X1 i_30_21 (.A1(n_30_13), .A2(n_30_14), .A3(n_30_15), .A4(n_30_16), 
      .ZN(n_309));
   NAND2_X1 i_30_22 (.A1(n_303), .A2(multiplicand[5]), .ZN(n_30_17));
   NAND2_X1 i_30_23 (.A1(n_301), .A2(n_52), .ZN(n_30_18));
   NAND2_X1 i_30_24 (.A1(n_302), .A2(n_51), .ZN(n_30_19));
   NAND2_X1 i_30_25 (.A1(n_304), .A2(multiplicand[4]), .ZN(n_30_20));
   NAND4_X1 i_30_26 (.A1(n_30_17), .A2(n_30_18), .A3(n_30_19), .A4(n_30_20), 
      .ZN(n_310));
   NAND2_X1 i_30_27 (.A1(n_303), .A2(multiplicand[6]), .ZN(n_30_21));
   NAND2_X1 i_30_28 (.A1(n_301), .A2(n_53), .ZN(n_30_22));
   NAND2_X1 i_30_29 (.A1(n_302), .A2(n_52), .ZN(n_30_23));
   NAND2_X1 i_30_30 (.A1(n_304), .A2(multiplicand[5]), .ZN(n_30_24));
   NAND4_X1 i_30_31 (.A1(n_30_21), .A2(n_30_22), .A3(n_30_23), .A4(n_30_24), 
      .ZN(n_311));
   NAND2_X1 i_30_32 (.A1(n_303), .A2(multiplicand[7]), .ZN(n_30_25));
   NAND2_X1 i_30_33 (.A1(n_301), .A2(n_54), .ZN(n_30_26));
   NAND2_X1 i_30_34 (.A1(n_302), .A2(n_53), .ZN(n_30_27));
   NAND2_X1 i_30_35 (.A1(n_304), .A2(multiplicand[6]), .ZN(n_30_28));
   NAND4_X1 i_30_36 (.A1(n_30_25), .A2(n_30_26), .A3(n_30_27), .A4(n_30_28), 
      .ZN(n_312));
   NAND2_X1 i_30_37 (.A1(n_303), .A2(multiplicand[8]), .ZN(n_30_29));
   NAND2_X1 i_30_38 (.A1(n_301), .A2(n_55), .ZN(n_30_30));
   NAND2_X1 i_30_39 (.A1(n_302), .A2(n_54), .ZN(n_30_31));
   NAND2_X1 i_30_40 (.A1(n_304), .A2(multiplicand[7]), .ZN(n_30_32));
   NAND4_X1 i_30_41 (.A1(n_30_29), .A2(n_30_30), .A3(n_30_31), .A4(n_30_32), 
      .ZN(n_313));
   NAND2_X1 i_30_42 (.A1(n_303), .A2(multiplicand[9]), .ZN(n_30_33));
   NAND2_X1 i_30_43 (.A1(n_301), .A2(n_56), .ZN(n_30_34));
   NAND2_X1 i_30_44 (.A1(n_302), .A2(n_55), .ZN(n_30_35));
   NAND2_X1 i_30_45 (.A1(n_304), .A2(multiplicand[8]), .ZN(n_30_36));
   NAND4_X1 i_30_46 (.A1(n_30_33), .A2(n_30_34), .A3(n_30_35), .A4(n_30_36), 
      .ZN(n_314));
   NAND2_X1 i_30_47 (.A1(n_303), .A2(multiplicand[10]), .ZN(n_30_37));
   NAND2_X1 i_30_48 (.A1(n_301), .A2(n_57), .ZN(n_30_38));
   NAND2_X1 i_30_49 (.A1(n_302), .A2(n_56), .ZN(n_30_39));
   NAND2_X1 i_30_50 (.A1(n_304), .A2(multiplicand[9]), .ZN(n_30_40));
   NAND4_X1 i_30_51 (.A1(n_30_37), .A2(n_30_38), .A3(n_30_39), .A4(n_30_40), 
      .ZN(n_315));
   NAND2_X1 i_30_52 (.A1(n_303), .A2(multiplicand[11]), .ZN(n_30_41));
   NAND2_X1 i_30_53 (.A1(n_301), .A2(n_58), .ZN(n_30_42));
   NAND2_X1 i_30_54 (.A1(n_302), .A2(n_57), .ZN(n_30_43));
   NAND2_X1 i_30_55 (.A1(n_304), .A2(multiplicand[10]), .ZN(n_30_44));
   NAND4_X1 i_30_56 (.A1(n_30_41), .A2(n_30_42), .A3(n_30_43), .A4(n_30_44), 
      .ZN(n_316));
   NAND2_X1 i_30_57 (.A1(n_303), .A2(multiplicand[12]), .ZN(n_30_45));
   NAND2_X1 i_30_58 (.A1(n_301), .A2(n_59), .ZN(n_30_46));
   NAND2_X1 i_30_59 (.A1(n_302), .A2(n_58), .ZN(n_30_47));
   NAND2_X1 i_30_60 (.A1(n_304), .A2(multiplicand[11]), .ZN(n_30_48));
   NAND4_X1 i_30_61 (.A1(n_30_45), .A2(n_30_46), .A3(n_30_47), .A4(n_30_48), 
      .ZN(n_317));
   NAND2_X1 i_30_62 (.A1(n_303), .A2(multiplicand[13]), .ZN(n_30_49));
   NAND2_X1 i_30_63 (.A1(n_301), .A2(n_60), .ZN(n_30_50));
   NAND2_X1 i_30_64 (.A1(n_302), .A2(n_59), .ZN(n_30_51));
   NAND2_X1 i_30_65 (.A1(n_304), .A2(multiplicand[12]), .ZN(n_30_52));
   NAND4_X1 i_30_66 (.A1(n_30_49), .A2(n_30_50), .A3(n_30_51), .A4(n_30_52), 
      .ZN(n_318));
   NAND2_X1 i_30_67 (.A1(n_303), .A2(multiplicand[14]), .ZN(n_30_53));
   NAND2_X1 i_30_68 (.A1(n_301), .A2(n_61), .ZN(n_30_54));
   NAND2_X1 i_30_69 (.A1(n_302), .A2(n_60), .ZN(n_30_55));
   NAND2_X1 i_30_70 (.A1(n_304), .A2(multiplicand[13]), .ZN(n_30_56));
   NAND4_X1 i_30_71 (.A1(n_30_53), .A2(n_30_54), .A3(n_30_55), .A4(n_30_56), 
      .ZN(n_319));
   NAND2_X1 i_30_72 (.A1(n_303), .A2(multiplicand[15]), .ZN(n_30_57));
   NAND2_X1 i_30_73 (.A1(n_301), .A2(n_62), .ZN(n_30_58));
   NAND2_X1 i_30_74 (.A1(n_302), .A2(n_61), .ZN(n_30_59));
   NAND2_X1 i_30_75 (.A1(n_304), .A2(multiplicand[14]), .ZN(n_30_60));
   NAND4_X1 i_30_76 (.A1(n_30_57), .A2(n_30_58), .A3(n_30_59), .A4(n_30_60), 
      .ZN(n_320));
   NAND2_X1 i_30_77 (.A1(n_303), .A2(multiplicand[16]), .ZN(n_30_61));
   NAND2_X1 i_30_78 (.A1(n_301), .A2(n_63), .ZN(n_30_62));
   NAND2_X1 i_30_79 (.A1(n_302), .A2(n_62), .ZN(n_30_63));
   NAND2_X1 i_30_80 (.A1(n_304), .A2(multiplicand[15]), .ZN(n_30_64));
   NAND4_X1 i_30_81 (.A1(n_30_61), .A2(n_30_62), .A3(n_30_63), .A4(n_30_64), 
      .ZN(n_321));
   NAND2_X1 i_30_82 (.A1(n_303), .A2(multiplicand[17]), .ZN(n_30_65));
   NAND2_X1 i_30_83 (.A1(n_301), .A2(n_64), .ZN(n_30_66));
   NAND2_X1 i_30_84 (.A1(n_302), .A2(n_63), .ZN(n_30_67));
   NAND2_X1 i_30_85 (.A1(n_304), .A2(multiplicand[16]), .ZN(n_30_68));
   NAND4_X1 i_30_86 (.A1(n_30_65), .A2(n_30_66), .A3(n_30_67), .A4(n_30_68), 
      .ZN(n_322));
   NAND2_X1 i_30_87 (.A1(n_303), .A2(multiplicand[18]), .ZN(n_30_69));
   NAND2_X1 i_30_88 (.A1(n_301), .A2(n_65), .ZN(n_30_70));
   NAND2_X1 i_30_89 (.A1(n_302), .A2(n_64), .ZN(n_30_71));
   NAND2_X1 i_30_90 (.A1(n_304), .A2(multiplicand[17]), .ZN(n_30_72));
   NAND4_X1 i_30_91 (.A1(n_30_69), .A2(n_30_70), .A3(n_30_71), .A4(n_30_72), 
      .ZN(n_323));
   NAND2_X1 i_30_92 (.A1(n_303), .A2(multiplicand[19]), .ZN(n_30_73));
   NAND2_X1 i_30_93 (.A1(n_301), .A2(n_66), .ZN(n_30_74));
   NAND2_X1 i_30_94 (.A1(n_302), .A2(n_65), .ZN(n_30_75));
   NAND2_X1 i_30_95 (.A1(n_304), .A2(multiplicand[18]), .ZN(n_30_76));
   NAND4_X1 i_30_96 (.A1(n_30_73), .A2(n_30_74), .A3(n_30_75), .A4(n_30_76), 
      .ZN(n_324));
   NAND2_X1 i_30_97 (.A1(n_303), .A2(multiplicand[20]), .ZN(n_30_77));
   NAND2_X1 i_30_98 (.A1(n_301), .A2(n_67), .ZN(n_30_78));
   NAND2_X1 i_30_99 (.A1(n_302), .A2(n_66), .ZN(n_30_79));
   NAND2_X1 i_30_100 (.A1(n_304), .A2(multiplicand[19]), .ZN(n_30_80));
   NAND4_X1 i_30_101 (.A1(n_30_77), .A2(n_30_78), .A3(n_30_79), .A4(n_30_80), 
      .ZN(n_325));
   NAND2_X1 i_30_102 (.A1(n_303), .A2(multiplicand[21]), .ZN(n_30_81));
   NAND2_X1 i_30_103 (.A1(n_301), .A2(n_68), .ZN(n_30_82));
   NAND2_X1 i_30_104 (.A1(n_302), .A2(n_67), .ZN(n_30_83));
   NAND2_X1 i_30_105 (.A1(n_304), .A2(multiplicand[20]), .ZN(n_30_84));
   NAND4_X1 i_30_106 (.A1(n_30_81), .A2(n_30_82), .A3(n_30_83), .A4(n_30_84), 
      .ZN(n_326));
   NAND2_X1 i_30_107 (.A1(n_303), .A2(multiplicand[22]), .ZN(n_30_85));
   NAND2_X1 i_30_108 (.A1(n_301), .A2(n_69), .ZN(n_30_86));
   NAND2_X1 i_30_109 (.A1(n_302), .A2(n_68), .ZN(n_30_87));
   NAND2_X1 i_30_110 (.A1(n_304), .A2(multiplicand[21]), .ZN(n_30_88));
   NAND4_X1 i_30_111 (.A1(n_30_85), .A2(n_30_86), .A3(n_30_87), .A4(n_30_88), 
      .ZN(n_327));
   NAND2_X1 i_30_112 (.A1(n_303), .A2(multiplicand[23]), .ZN(n_30_89));
   NAND2_X1 i_30_113 (.A1(n_301), .A2(n_70), .ZN(n_30_90));
   NAND2_X1 i_30_114 (.A1(n_302), .A2(n_69), .ZN(n_30_91));
   NAND2_X1 i_30_115 (.A1(n_304), .A2(multiplicand[22]), .ZN(n_30_92));
   NAND4_X1 i_30_116 (.A1(n_30_89), .A2(n_30_90), .A3(n_30_91), .A4(n_30_92), 
      .ZN(n_328));
   NAND2_X1 i_30_117 (.A1(n_303), .A2(multiplicand[24]), .ZN(n_30_93));
   NAND2_X1 i_30_118 (.A1(n_301), .A2(n_71), .ZN(n_30_94));
   NAND2_X1 i_30_119 (.A1(n_302), .A2(n_70), .ZN(n_30_95));
   NAND2_X1 i_30_120 (.A1(n_304), .A2(multiplicand[23]), .ZN(n_30_96));
   NAND4_X1 i_30_121 (.A1(n_30_93), .A2(n_30_94), .A3(n_30_95), .A4(n_30_96), 
      .ZN(n_329));
   NAND2_X1 i_30_122 (.A1(n_303), .A2(multiplicand[25]), .ZN(n_30_97));
   NAND2_X1 i_30_123 (.A1(n_301), .A2(n_72), .ZN(n_30_98));
   NAND2_X1 i_30_124 (.A1(n_302), .A2(n_71), .ZN(n_30_99));
   NAND2_X1 i_30_125 (.A1(n_304), .A2(multiplicand[24]), .ZN(n_30_100));
   NAND4_X1 i_30_126 (.A1(n_30_97), .A2(n_30_98), .A3(n_30_99), .A4(n_30_100), 
      .ZN(n_330));
   NAND2_X1 i_30_127 (.A1(n_303), .A2(multiplicand[26]), .ZN(n_30_101));
   NAND2_X1 i_30_128 (.A1(n_301), .A2(n_73), .ZN(n_30_102));
   NAND2_X1 i_30_129 (.A1(n_302), .A2(n_72), .ZN(n_30_103));
   NAND2_X1 i_30_130 (.A1(n_304), .A2(multiplicand[25]), .ZN(n_30_104));
   NAND4_X1 i_30_131 (.A1(n_30_101), .A2(n_30_102), .A3(n_30_103), .A4(n_30_104), 
      .ZN(n_331));
   NAND2_X1 i_30_132 (.A1(n_303), .A2(multiplicand[27]), .ZN(n_30_105));
   NAND2_X1 i_30_133 (.A1(n_301), .A2(n_74), .ZN(n_30_106));
   NAND2_X1 i_30_134 (.A1(n_302), .A2(n_73), .ZN(n_30_107));
   NAND2_X1 i_30_135 (.A1(n_304), .A2(multiplicand[26]), .ZN(n_30_108));
   NAND4_X1 i_30_136 (.A1(n_30_105), .A2(n_30_106), .A3(n_30_107), .A4(n_30_108), 
      .ZN(n_332));
   NAND2_X1 i_30_137 (.A1(n_303), .A2(multiplicand[28]), .ZN(n_30_109));
   NAND2_X1 i_30_138 (.A1(n_301), .A2(n_75), .ZN(n_30_110));
   NAND2_X1 i_30_139 (.A1(n_302), .A2(n_74), .ZN(n_30_111));
   NAND2_X1 i_30_140 (.A1(n_304), .A2(multiplicand[27]), .ZN(n_30_112));
   NAND4_X1 i_30_141 (.A1(n_30_109), .A2(n_30_110), .A3(n_30_111), .A4(n_30_112), 
      .ZN(n_333));
   NAND2_X1 i_30_142 (.A1(n_303), .A2(multiplicand[29]), .ZN(n_30_113));
   NAND2_X1 i_30_143 (.A1(n_301), .A2(n_76), .ZN(n_30_114));
   NAND2_X1 i_30_144 (.A1(n_302), .A2(n_75), .ZN(n_30_115));
   NAND2_X1 i_30_145 (.A1(n_304), .A2(multiplicand[28]), .ZN(n_30_116));
   NAND4_X1 i_30_146 (.A1(n_30_113), .A2(n_30_114), .A3(n_30_115), .A4(n_30_116), 
      .ZN(n_334));
   NAND2_X1 i_30_147 (.A1(n_303), .A2(multiplicand[30]), .ZN(n_30_117));
   NAND2_X1 i_30_148 (.A1(n_301), .A2(n_77), .ZN(n_30_118));
   NAND2_X1 i_30_149 (.A1(n_302), .A2(n_76), .ZN(n_30_119));
   NAND2_X1 i_30_150 (.A1(n_304), .A2(multiplicand[29]), .ZN(n_30_120));
   NAND4_X1 i_30_151 (.A1(n_30_117), .A2(n_30_118), .A3(n_30_119), .A4(n_30_120), 
      .ZN(n_335));
   NAND2_X1 i_30_152 (.A1(n_303), .A2(multiplicand[31]), .ZN(n_30_121));
   NAND2_X1 i_30_153 (.A1(n_301), .A2(n_78), .ZN(n_30_122));
   NAND2_X1 i_30_154 (.A1(n_302), .A2(n_77), .ZN(n_30_123));
   NAND2_X1 i_30_155 (.A1(n_304), .A2(multiplicand[30]), .ZN(n_30_124));
   NAND4_X1 i_30_156 (.A1(n_30_121), .A2(n_30_122), .A3(n_30_123), .A4(n_30_124), 
      .ZN(n_336));
   NAND2_X1 i_30_157 (.A1(n_302), .A2(n_78), .ZN(n_30_125));
   NAND2_X1 i_30_158 (.A1(n_304), .A2(multiplicand[31]), .ZN(n_30_126));
   NAND4_X1 i_30_159 (.A1(n_30_121), .A2(n_30_122), .A3(n_30_125), .A4(n_30_126), 
      .ZN(n_337));
   INV_X1 i_31_0 (.A(n_21), .ZN(n_31_0));
   AND3_X1 i_31_1 (.A1(n_31_0), .A2(n_22), .A3(n_23), .ZN(n_338));
   INV_X1 i_31_2 (.A(n_22), .ZN(n_31_1));
   AND3_X1 i_31_3 (.A1(n_31_1), .A2(n_21), .A3(n_23), .ZN(n_339));
   NOR3_X1 i_31_4 (.A1(n_31_1), .A2(n_21), .A3(n_23), .ZN(n_340));
   NOR3_X1 i_31_5 (.A1(n_31_0), .A2(n_22), .A3(n_23), .ZN(n_341));
   AOI22_X1 i_32_0 (.A1(n_340), .A2(multiplicand[0]), .B1(n_338), .B2(
      multiplicand[0]), .ZN(n_32_0));
   INV_X1 i_32_1 (.A(n_32_0), .ZN(n_342));
   NAND2_X1 i_32_2 (.A1(n_340), .A2(multiplicand[1]), .ZN(n_32_1));
   NAND2_X1 i_32_3 (.A1(n_338), .A2(n_48), .ZN(n_32_2));
   NAND2_X1 i_32_4 (.A1(n_339), .A2(multiplicand[0]), .ZN(n_32_3));
   NAND2_X1 i_32_5 (.A1(n_341), .A2(multiplicand[0]), .ZN(n_32_4));
   NAND4_X1 i_32_6 (.A1(n_32_1), .A2(n_32_2), .A3(n_32_3), .A4(n_32_4), .ZN(
      n_343));
   NAND2_X1 i_32_7 (.A1(n_340), .A2(multiplicand[2]), .ZN(n_32_5));
   NAND2_X1 i_32_8 (.A1(n_338), .A2(n_49), .ZN(n_32_6));
   NAND2_X1 i_32_9 (.A1(n_339), .A2(n_48), .ZN(n_32_7));
   NAND2_X1 i_32_10 (.A1(n_341), .A2(multiplicand[1]), .ZN(n_32_8));
   NAND4_X1 i_32_11 (.A1(n_32_5), .A2(n_32_6), .A3(n_32_7), .A4(n_32_8), 
      .ZN(n_344));
   NAND2_X1 i_32_12 (.A1(n_340), .A2(multiplicand[3]), .ZN(n_32_9));
   NAND2_X1 i_32_13 (.A1(n_338), .A2(n_50), .ZN(n_32_10));
   NAND2_X1 i_32_14 (.A1(n_339), .A2(n_49), .ZN(n_32_11));
   NAND2_X1 i_32_15 (.A1(n_341), .A2(multiplicand[2]), .ZN(n_32_12));
   NAND4_X1 i_32_16 (.A1(n_32_9), .A2(n_32_10), .A3(n_32_11), .A4(n_32_12), 
      .ZN(n_345));
   NAND2_X1 i_32_17 (.A1(n_340), .A2(multiplicand[4]), .ZN(n_32_13));
   NAND2_X1 i_32_18 (.A1(n_338), .A2(n_51), .ZN(n_32_14));
   NAND2_X1 i_32_19 (.A1(n_339), .A2(n_50), .ZN(n_32_15));
   NAND2_X1 i_32_20 (.A1(n_341), .A2(multiplicand[3]), .ZN(n_32_16));
   NAND4_X1 i_32_21 (.A1(n_32_13), .A2(n_32_14), .A3(n_32_15), .A4(n_32_16), 
      .ZN(n_346));
   NAND2_X1 i_32_22 (.A1(n_340), .A2(multiplicand[5]), .ZN(n_32_17));
   NAND2_X1 i_32_23 (.A1(n_338), .A2(n_52), .ZN(n_32_18));
   NAND2_X1 i_32_24 (.A1(n_339), .A2(n_51), .ZN(n_32_19));
   NAND2_X1 i_32_25 (.A1(n_341), .A2(multiplicand[4]), .ZN(n_32_20));
   NAND4_X1 i_32_26 (.A1(n_32_17), .A2(n_32_18), .A3(n_32_19), .A4(n_32_20), 
      .ZN(n_347));
   NAND2_X1 i_32_27 (.A1(n_340), .A2(multiplicand[6]), .ZN(n_32_21));
   NAND2_X1 i_32_28 (.A1(n_338), .A2(n_53), .ZN(n_32_22));
   NAND2_X1 i_32_29 (.A1(n_339), .A2(n_52), .ZN(n_32_23));
   NAND2_X1 i_32_30 (.A1(n_341), .A2(multiplicand[5]), .ZN(n_32_24));
   NAND4_X1 i_32_31 (.A1(n_32_21), .A2(n_32_22), .A3(n_32_23), .A4(n_32_24), 
      .ZN(n_348));
   NAND2_X1 i_32_32 (.A1(n_340), .A2(multiplicand[7]), .ZN(n_32_25));
   NAND2_X1 i_32_33 (.A1(n_338), .A2(n_54), .ZN(n_32_26));
   NAND2_X1 i_32_34 (.A1(n_339), .A2(n_53), .ZN(n_32_27));
   NAND2_X1 i_32_35 (.A1(n_341), .A2(multiplicand[6]), .ZN(n_32_28));
   NAND4_X1 i_32_36 (.A1(n_32_25), .A2(n_32_26), .A3(n_32_27), .A4(n_32_28), 
      .ZN(n_349));
   NAND2_X1 i_32_37 (.A1(n_340), .A2(multiplicand[8]), .ZN(n_32_29));
   NAND2_X1 i_32_38 (.A1(n_338), .A2(n_55), .ZN(n_32_30));
   NAND2_X1 i_32_39 (.A1(n_339), .A2(n_54), .ZN(n_32_31));
   NAND2_X1 i_32_40 (.A1(n_341), .A2(multiplicand[7]), .ZN(n_32_32));
   NAND4_X1 i_32_41 (.A1(n_32_29), .A2(n_32_30), .A3(n_32_31), .A4(n_32_32), 
      .ZN(n_350));
   NAND2_X1 i_32_42 (.A1(n_340), .A2(multiplicand[9]), .ZN(n_32_33));
   NAND2_X1 i_32_43 (.A1(n_338), .A2(n_56), .ZN(n_32_34));
   NAND2_X1 i_32_44 (.A1(n_339), .A2(n_55), .ZN(n_32_35));
   NAND2_X1 i_32_45 (.A1(n_341), .A2(multiplicand[8]), .ZN(n_32_36));
   NAND4_X1 i_32_46 (.A1(n_32_33), .A2(n_32_34), .A3(n_32_35), .A4(n_32_36), 
      .ZN(n_351));
   NAND2_X1 i_32_47 (.A1(n_340), .A2(multiplicand[10]), .ZN(n_32_37));
   NAND2_X1 i_32_48 (.A1(n_338), .A2(n_57), .ZN(n_32_38));
   NAND2_X1 i_32_49 (.A1(n_339), .A2(n_56), .ZN(n_32_39));
   NAND2_X1 i_32_50 (.A1(n_341), .A2(multiplicand[9]), .ZN(n_32_40));
   NAND4_X1 i_32_51 (.A1(n_32_37), .A2(n_32_38), .A3(n_32_39), .A4(n_32_40), 
      .ZN(n_352));
   NAND2_X1 i_32_52 (.A1(n_340), .A2(multiplicand[11]), .ZN(n_32_41));
   NAND2_X1 i_32_53 (.A1(n_338), .A2(n_58), .ZN(n_32_42));
   NAND2_X1 i_32_54 (.A1(n_339), .A2(n_57), .ZN(n_32_43));
   NAND2_X1 i_32_55 (.A1(n_341), .A2(multiplicand[10]), .ZN(n_32_44));
   NAND4_X1 i_32_56 (.A1(n_32_41), .A2(n_32_42), .A3(n_32_43), .A4(n_32_44), 
      .ZN(n_353));
   NAND2_X1 i_32_57 (.A1(n_340), .A2(multiplicand[12]), .ZN(n_32_45));
   NAND2_X1 i_32_58 (.A1(n_338), .A2(n_59), .ZN(n_32_46));
   NAND2_X1 i_32_59 (.A1(n_339), .A2(n_58), .ZN(n_32_47));
   NAND2_X1 i_32_60 (.A1(n_341), .A2(multiplicand[11]), .ZN(n_32_48));
   NAND4_X1 i_32_61 (.A1(n_32_45), .A2(n_32_46), .A3(n_32_47), .A4(n_32_48), 
      .ZN(n_354));
   NAND2_X1 i_32_62 (.A1(n_340), .A2(multiplicand[13]), .ZN(n_32_49));
   NAND2_X1 i_32_63 (.A1(n_338), .A2(n_60), .ZN(n_32_50));
   NAND2_X1 i_32_64 (.A1(n_339), .A2(n_59), .ZN(n_32_51));
   NAND2_X1 i_32_65 (.A1(n_341), .A2(multiplicand[12]), .ZN(n_32_52));
   NAND4_X1 i_32_66 (.A1(n_32_49), .A2(n_32_50), .A3(n_32_51), .A4(n_32_52), 
      .ZN(n_355));
   NAND2_X1 i_32_67 (.A1(n_340), .A2(multiplicand[14]), .ZN(n_32_53));
   NAND2_X1 i_32_68 (.A1(n_338), .A2(n_61), .ZN(n_32_54));
   NAND2_X1 i_32_69 (.A1(n_339), .A2(n_60), .ZN(n_32_55));
   NAND2_X1 i_32_70 (.A1(n_341), .A2(multiplicand[13]), .ZN(n_32_56));
   NAND4_X1 i_32_71 (.A1(n_32_53), .A2(n_32_54), .A3(n_32_55), .A4(n_32_56), 
      .ZN(n_356));
   NAND2_X1 i_32_72 (.A1(n_340), .A2(multiplicand[15]), .ZN(n_32_57));
   NAND2_X1 i_32_73 (.A1(n_338), .A2(n_62), .ZN(n_32_58));
   NAND2_X1 i_32_74 (.A1(n_339), .A2(n_61), .ZN(n_32_59));
   NAND2_X1 i_32_75 (.A1(n_341), .A2(multiplicand[14]), .ZN(n_32_60));
   NAND4_X1 i_32_76 (.A1(n_32_57), .A2(n_32_58), .A3(n_32_59), .A4(n_32_60), 
      .ZN(n_357));
   NAND2_X1 i_32_77 (.A1(n_340), .A2(multiplicand[16]), .ZN(n_32_61));
   NAND2_X1 i_32_78 (.A1(n_338), .A2(n_63), .ZN(n_32_62));
   NAND2_X1 i_32_79 (.A1(n_339), .A2(n_62), .ZN(n_32_63));
   NAND2_X1 i_32_80 (.A1(n_341), .A2(multiplicand[15]), .ZN(n_32_64));
   NAND4_X1 i_32_81 (.A1(n_32_61), .A2(n_32_62), .A3(n_32_63), .A4(n_32_64), 
      .ZN(n_358));
   NAND2_X1 i_32_82 (.A1(n_340), .A2(multiplicand[17]), .ZN(n_32_65));
   NAND2_X1 i_32_83 (.A1(n_338), .A2(n_64), .ZN(n_32_66));
   NAND2_X1 i_32_84 (.A1(n_339), .A2(n_63), .ZN(n_32_67));
   NAND2_X1 i_32_85 (.A1(n_341), .A2(multiplicand[16]), .ZN(n_32_68));
   NAND4_X1 i_32_86 (.A1(n_32_65), .A2(n_32_66), .A3(n_32_67), .A4(n_32_68), 
      .ZN(n_359));
   NAND2_X1 i_32_87 (.A1(n_340), .A2(multiplicand[18]), .ZN(n_32_69));
   NAND2_X1 i_32_88 (.A1(n_338), .A2(n_65), .ZN(n_32_70));
   NAND2_X1 i_32_89 (.A1(n_339), .A2(n_64), .ZN(n_32_71));
   NAND2_X1 i_32_90 (.A1(n_341), .A2(multiplicand[17]), .ZN(n_32_72));
   NAND4_X1 i_32_91 (.A1(n_32_69), .A2(n_32_70), .A3(n_32_71), .A4(n_32_72), 
      .ZN(n_360));
   NAND2_X1 i_32_92 (.A1(n_340), .A2(multiplicand[19]), .ZN(n_32_73));
   NAND2_X1 i_32_93 (.A1(n_338), .A2(n_66), .ZN(n_32_74));
   NAND2_X1 i_32_94 (.A1(n_339), .A2(n_65), .ZN(n_32_75));
   NAND2_X1 i_32_95 (.A1(n_341), .A2(multiplicand[18]), .ZN(n_32_76));
   NAND4_X1 i_32_96 (.A1(n_32_73), .A2(n_32_74), .A3(n_32_75), .A4(n_32_76), 
      .ZN(n_361));
   NAND2_X1 i_32_97 (.A1(n_340), .A2(multiplicand[20]), .ZN(n_32_77));
   NAND2_X1 i_32_98 (.A1(n_338), .A2(n_67), .ZN(n_32_78));
   NAND2_X1 i_32_99 (.A1(n_339), .A2(n_66), .ZN(n_32_79));
   NAND2_X1 i_32_100 (.A1(n_341), .A2(multiplicand[19]), .ZN(n_32_80));
   NAND4_X1 i_32_101 (.A1(n_32_77), .A2(n_32_78), .A3(n_32_79), .A4(n_32_80), 
      .ZN(n_362));
   NAND2_X1 i_32_102 (.A1(n_340), .A2(multiplicand[21]), .ZN(n_32_81));
   NAND2_X1 i_32_103 (.A1(n_338), .A2(n_68), .ZN(n_32_82));
   NAND2_X1 i_32_104 (.A1(n_339), .A2(n_67), .ZN(n_32_83));
   NAND2_X1 i_32_105 (.A1(n_341), .A2(multiplicand[20]), .ZN(n_32_84));
   NAND4_X1 i_32_106 (.A1(n_32_81), .A2(n_32_82), .A3(n_32_83), .A4(n_32_84), 
      .ZN(n_363));
   NAND2_X1 i_32_107 (.A1(n_340), .A2(multiplicand[22]), .ZN(n_32_85));
   NAND2_X1 i_32_108 (.A1(n_338), .A2(n_69), .ZN(n_32_86));
   NAND2_X1 i_32_109 (.A1(n_339), .A2(n_68), .ZN(n_32_87));
   NAND2_X1 i_32_110 (.A1(n_341), .A2(multiplicand[21]), .ZN(n_32_88));
   NAND4_X1 i_32_111 (.A1(n_32_85), .A2(n_32_86), .A3(n_32_87), .A4(n_32_88), 
      .ZN(n_364));
   NAND2_X1 i_32_112 (.A1(n_340), .A2(multiplicand[23]), .ZN(n_32_89));
   NAND2_X1 i_32_113 (.A1(n_338), .A2(n_70), .ZN(n_32_90));
   NAND2_X1 i_32_114 (.A1(n_339), .A2(n_69), .ZN(n_32_91));
   NAND2_X1 i_32_115 (.A1(n_341), .A2(multiplicand[22]), .ZN(n_32_92));
   NAND4_X1 i_32_116 (.A1(n_32_89), .A2(n_32_90), .A3(n_32_91), .A4(n_32_92), 
      .ZN(n_365));
   NAND2_X1 i_32_117 (.A1(n_340), .A2(multiplicand[24]), .ZN(n_32_93));
   NAND2_X1 i_32_118 (.A1(n_338), .A2(n_71), .ZN(n_32_94));
   NAND2_X1 i_32_119 (.A1(n_339), .A2(n_70), .ZN(n_32_95));
   NAND2_X1 i_32_120 (.A1(n_341), .A2(multiplicand[23]), .ZN(n_32_96));
   NAND4_X1 i_32_121 (.A1(n_32_93), .A2(n_32_94), .A3(n_32_95), .A4(n_32_96), 
      .ZN(n_366));
   NAND2_X1 i_32_122 (.A1(n_340), .A2(multiplicand[25]), .ZN(n_32_97));
   NAND2_X1 i_32_123 (.A1(n_338), .A2(n_72), .ZN(n_32_98));
   NAND2_X1 i_32_124 (.A1(n_339), .A2(n_71), .ZN(n_32_99));
   NAND2_X1 i_32_125 (.A1(n_341), .A2(multiplicand[24]), .ZN(n_32_100));
   NAND4_X1 i_32_126 (.A1(n_32_97), .A2(n_32_98), .A3(n_32_99), .A4(n_32_100), 
      .ZN(n_367));
   NAND2_X1 i_32_127 (.A1(n_340), .A2(multiplicand[26]), .ZN(n_32_101));
   NAND2_X1 i_32_128 (.A1(n_338), .A2(n_73), .ZN(n_32_102));
   NAND2_X1 i_32_129 (.A1(n_339), .A2(n_72), .ZN(n_32_103));
   NAND2_X1 i_32_130 (.A1(n_341), .A2(multiplicand[25]), .ZN(n_32_104));
   NAND4_X1 i_32_131 (.A1(n_32_101), .A2(n_32_102), .A3(n_32_103), .A4(n_32_104), 
      .ZN(n_368));
   NAND2_X1 i_32_132 (.A1(n_340), .A2(multiplicand[27]), .ZN(n_32_105));
   NAND2_X1 i_32_133 (.A1(n_338), .A2(n_74), .ZN(n_32_106));
   NAND2_X1 i_32_134 (.A1(n_339), .A2(n_73), .ZN(n_32_107));
   NAND2_X1 i_32_135 (.A1(n_341), .A2(multiplicand[26]), .ZN(n_32_108));
   NAND4_X1 i_32_136 (.A1(n_32_105), .A2(n_32_106), .A3(n_32_107), .A4(n_32_108), 
      .ZN(n_369));
   NAND2_X1 i_32_137 (.A1(n_340), .A2(multiplicand[28]), .ZN(n_32_109));
   NAND2_X1 i_32_138 (.A1(n_338), .A2(n_75), .ZN(n_32_110));
   NAND2_X1 i_32_139 (.A1(n_339), .A2(n_74), .ZN(n_32_111));
   NAND2_X1 i_32_140 (.A1(n_341), .A2(multiplicand[27]), .ZN(n_32_112));
   NAND4_X1 i_32_141 (.A1(n_32_109), .A2(n_32_110), .A3(n_32_111), .A4(n_32_112), 
      .ZN(n_370));
   NAND2_X1 i_32_142 (.A1(n_340), .A2(multiplicand[29]), .ZN(n_32_113));
   NAND2_X1 i_32_143 (.A1(n_338), .A2(n_76), .ZN(n_32_114));
   NAND2_X1 i_32_144 (.A1(n_339), .A2(n_75), .ZN(n_32_115));
   NAND2_X1 i_32_145 (.A1(n_341), .A2(multiplicand[28]), .ZN(n_32_116));
   NAND4_X1 i_32_146 (.A1(n_32_113), .A2(n_32_114), .A3(n_32_115), .A4(n_32_116), 
      .ZN(n_371));
   NAND2_X1 i_32_147 (.A1(n_340), .A2(multiplicand[30]), .ZN(n_32_117));
   NAND2_X1 i_32_148 (.A1(n_338), .A2(n_77), .ZN(n_32_118));
   NAND2_X1 i_32_149 (.A1(n_339), .A2(n_76), .ZN(n_32_119));
   NAND2_X1 i_32_150 (.A1(n_341), .A2(multiplicand[29]), .ZN(n_32_120));
   NAND4_X1 i_32_151 (.A1(n_32_117), .A2(n_32_118), .A3(n_32_119), .A4(n_32_120), 
      .ZN(n_372));
   NAND2_X1 i_32_152 (.A1(n_340), .A2(multiplicand[31]), .ZN(n_32_121));
   NAND2_X1 i_32_153 (.A1(n_338), .A2(n_78), .ZN(n_32_122));
   NAND2_X1 i_32_154 (.A1(n_339), .A2(n_77), .ZN(n_32_123));
   NAND2_X1 i_32_155 (.A1(n_341), .A2(multiplicand[30]), .ZN(n_32_124));
   NAND4_X1 i_32_156 (.A1(n_32_121), .A2(n_32_122), .A3(n_32_123), .A4(n_32_124), 
      .ZN(n_373));
   NAND2_X1 i_32_157 (.A1(n_339), .A2(n_78), .ZN(n_32_125));
   NAND2_X1 i_32_158 (.A1(n_341), .A2(multiplicand[31]), .ZN(n_32_126));
   NAND4_X1 i_32_159 (.A1(n_32_121), .A2(n_32_122), .A3(n_32_125), .A4(n_32_126), 
      .ZN(n_374));
   INV_X1 i_33_0 (.A(n_24), .ZN(n_33_0));
   AND3_X1 i_33_1 (.A1(n_33_0), .A2(n_25), .A3(n_26), .ZN(n_375));
   INV_X1 i_33_2 (.A(n_25), .ZN(n_33_1));
   AND3_X1 i_33_3 (.A1(n_33_1), .A2(n_24), .A3(n_26), .ZN(n_376));
   NOR3_X1 i_33_4 (.A1(n_33_1), .A2(n_24), .A3(n_26), .ZN(n_377));
   NOR3_X1 i_33_5 (.A1(n_33_0), .A2(n_25), .A3(n_26), .ZN(n_378));
   AOI22_X1 i_34_0 (.A1(n_377), .A2(multiplicand[0]), .B1(n_375), .B2(
      multiplicand[0]), .ZN(n_34_0));
   INV_X1 i_34_1 (.A(n_34_0), .ZN(n_379));
   NAND2_X1 i_34_2 (.A1(n_377), .A2(multiplicand[1]), .ZN(n_34_1));
   NAND2_X1 i_34_3 (.A1(n_375), .A2(n_48), .ZN(n_34_2));
   NAND2_X1 i_34_4 (.A1(n_376), .A2(multiplicand[0]), .ZN(n_34_3));
   NAND2_X1 i_34_5 (.A1(n_378), .A2(multiplicand[0]), .ZN(n_34_4));
   NAND4_X1 i_34_6 (.A1(n_34_1), .A2(n_34_2), .A3(n_34_3), .A4(n_34_4), .ZN(
      n_380));
   NAND2_X1 i_34_7 (.A1(n_377), .A2(multiplicand[2]), .ZN(n_34_5));
   NAND2_X1 i_34_8 (.A1(n_375), .A2(n_49), .ZN(n_34_6));
   NAND2_X1 i_34_9 (.A1(n_376), .A2(n_48), .ZN(n_34_7));
   NAND2_X1 i_34_10 (.A1(n_378), .A2(multiplicand[1]), .ZN(n_34_8));
   NAND4_X1 i_34_11 (.A1(n_34_5), .A2(n_34_6), .A3(n_34_7), .A4(n_34_8), 
      .ZN(n_381));
   NAND2_X1 i_34_12 (.A1(n_377), .A2(multiplicand[3]), .ZN(n_34_9));
   NAND2_X1 i_34_13 (.A1(n_375), .A2(n_50), .ZN(n_34_10));
   NAND2_X1 i_34_14 (.A1(n_376), .A2(n_49), .ZN(n_34_11));
   NAND2_X1 i_34_15 (.A1(n_378), .A2(multiplicand[2]), .ZN(n_34_12));
   NAND4_X1 i_34_16 (.A1(n_34_9), .A2(n_34_10), .A3(n_34_11), .A4(n_34_12), 
      .ZN(n_382));
   NAND2_X1 i_34_17 (.A1(n_377), .A2(multiplicand[4]), .ZN(n_34_13));
   NAND2_X1 i_34_18 (.A1(n_375), .A2(n_51), .ZN(n_34_14));
   NAND2_X1 i_34_19 (.A1(n_376), .A2(n_50), .ZN(n_34_15));
   NAND2_X1 i_34_20 (.A1(n_378), .A2(multiplicand[3]), .ZN(n_34_16));
   NAND4_X1 i_34_21 (.A1(n_34_13), .A2(n_34_14), .A3(n_34_15), .A4(n_34_16), 
      .ZN(n_383));
   NAND2_X1 i_34_22 (.A1(n_377), .A2(multiplicand[5]), .ZN(n_34_17));
   NAND2_X1 i_34_23 (.A1(n_375), .A2(n_52), .ZN(n_34_18));
   NAND2_X1 i_34_24 (.A1(n_376), .A2(n_51), .ZN(n_34_19));
   NAND2_X1 i_34_25 (.A1(n_378), .A2(multiplicand[4]), .ZN(n_34_20));
   NAND4_X1 i_34_26 (.A1(n_34_17), .A2(n_34_18), .A3(n_34_19), .A4(n_34_20), 
      .ZN(n_384));
   NAND2_X1 i_34_27 (.A1(n_377), .A2(multiplicand[6]), .ZN(n_34_21));
   NAND2_X1 i_34_28 (.A1(n_375), .A2(n_53), .ZN(n_34_22));
   NAND2_X1 i_34_29 (.A1(n_376), .A2(n_52), .ZN(n_34_23));
   NAND2_X1 i_34_30 (.A1(n_378), .A2(multiplicand[5]), .ZN(n_34_24));
   NAND4_X1 i_34_31 (.A1(n_34_21), .A2(n_34_22), .A3(n_34_23), .A4(n_34_24), 
      .ZN(n_385));
   NAND2_X1 i_34_32 (.A1(n_377), .A2(multiplicand[7]), .ZN(n_34_25));
   NAND2_X1 i_34_33 (.A1(n_375), .A2(n_54), .ZN(n_34_26));
   NAND2_X1 i_34_34 (.A1(n_376), .A2(n_53), .ZN(n_34_27));
   NAND2_X1 i_34_35 (.A1(n_378), .A2(multiplicand[6]), .ZN(n_34_28));
   NAND4_X1 i_34_36 (.A1(n_34_25), .A2(n_34_26), .A3(n_34_27), .A4(n_34_28), 
      .ZN(n_386));
   NAND2_X1 i_34_37 (.A1(n_377), .A2(multiplicand[8]), .ZN(n_34_29));
   NAND2_X1 i_34_38 (.A1(n_375), .A2(n_55), .ZN(n_34_30));
   NAND2_X1 i_34_39 (.A1(n_376), .A2(n_54), .ZN(n_34_31));
   NAND2_X1 i_34_40 (.A1(n_378), .A2(multiplicand[7]), .ZN(n_34_32));
   NAND4_X1 i_34_41 (.A1(n_34_29), .A2(n_34_30), .A3(n_34_31), .A4(n_34_32), 
      .ZN(n_387));
   NAND2_X1 i_34_42 (.A1(n_377), .A2(multiplicand[9]), .ZN(n_34_33));
   NAND2_X1 i_34_43 (.A1(n_375), .A2(n_56), .ZN(n_34_34));
   NAND2_X1 i_34_44 (.A1(n_376), .A2(n_55), .ZN(n_34_35));
   NAND2_X1 i_34_45 (.A1(n_378), .A2(multiplicand[8]), .ZN(n_34_36));
   NAND4_X1 i_34_46 (.A1(n_34_33), .A2(n_34_34), .A3(n_34_35), .A4(n_34_36), 
      .ZN(n_388));
   NAND2_X1 i_34_47 (.A1(n_377), .A2(multiplicand[10]), .ZN(n_34_37));
   NAND2_X1 i_34_48 (.A1(n_375), .A2(n_57), .ZN(n_34_38));
   NAND2_X1 i_34_49 (.A1(n_376), .A2(n_56), .ZN(n_34_39));
   NAND2_X1 i_34_50 (.A1(n_378), .A2(multiplicand[9]), .ZN(n_34_40));
   NAND4_X1 i_34_51 (.A1(n_34_37), .A2(n_34_38), .A3(n_34_39), .A4(n_34_40), 
      .ZN(n_389));
   NAND2_X1 i_34_52 (.A1(n_377), .A2(multiplicand[11]), .ZN(n_34_41));
   NAND2_X1 i_34_53 (.A1(n_375), .A2(n_58), .ZN(n_34_42));
   NAND2_X1 i_34_54 (.A1(n_376), .A2(n_57), .ZN(n_34_43));
   NAND2_X1 i_34_55 (.A1(n_378), .A2(multiplicand[10]), .ZN(n_34_44));
   NAND4_X1 i_34_56 (.A1(n_34_41), .A2(n_34_42), .A3(n_34_43), .A4(n_34_44), 
      .ZN(n_390));
   NAND2_X1 i_34_57 (.A1(n_377), .A2(multiplicand[12]), .ZN(n_34_45));
   NAND2_X1 i_34_58 (.A1(n_375), .A2(n_59), .ZN(n_34_46));
   NAND2_X1 i_34_59 (.A1(n_376), .A2(n_58), .ZN(n_34_47));
   NAND2_X1 i_34_60 (.A1(n_378), .A2(multiplicand[11]), .ZN(n_34_48));
   NAND4_X1 i_34_61 (.A1(n_34_45), .A2(n_34_46), .A3(n_34_47), .A4(n_34_48), 
      .ZN(n_391));
   NAND2_X1 i_34_62 (.A1(n_377), .A2(multiplicand[13]), .ZN(n_34_49));
   NAND2_X1 i_34_63 (.A1(n_375), .A2(n_60), .ZN(n_34_50));
   NAND2_X1 i_34_64 (.A1(n_376), .A2(n_59), .ZN(n_34_51));
   NAND2_X1 i_34_65 (.A1(n_378), .A2(multiplicand[12]), .ZN(n_34_52));
   NAND4_X1 i_34_66 (.A1(n_34_49), .A2(n_34_50), .A3(n_34_51), .A4(n_34_52), 
      .ZN(n_392));
   NAND2_X1 i_34_67 (.A1(n_377), .A2(multiplicand[14]), .ZN(n_34_53));
   NAND2_X1 i_34_68 (.A1(n_375), .A2(n_61), .ZN(n_34_54));
   NAND2_X1 i_34_69 (.A1(n_376), .A2(n_60), .ZN(n_34_55));
   NAND2_X1 i_34_70 (.A1(n_378), .A2(multiplicand[13]), .ZN(n_34_56));
   NAND4_X1 i_34_71 (.A1(n_34_53), .A2(n_34_54), .A3(n_34_55), .A4(n_34_56), 
      .ZN(n_393));
   NAND2_X1 i_34_72 (.A1(n_377), .A2(multiplicand[15]), .ZN(n_34_57));
   NAND2_X1 i_34_73 (.A1(n_375), .A2(n_62), .ZN(n_34_58));
   NAND2_X1 i_34_74 (.A1(n_376), .A2(n_61), .ZN(n_34_59));
   NAND2_X1 i_34_75 (.A1(n_378), .A2(multiplicand[14]), .ZN(n_34_60));
   NAND4_X1 i_34_76 (.A1(n_34_57), .A2(n_34_58), .A3(n_34_59), .A4(n_34_60), 
      .ZN(n_394));
   NAND2_X1 i_34_77 (.A1(n_377), .A2(multiplicand[16]), .ZN(n_34_61));
   NAND2_X1 i_34_78 (.A1(n_375), .A2(n_63), .ZN(n_34_62));
   NAND2_X1 i_34_79 (.A1(n_376), .A2(n_62), .ZN(n_34_63));
   NAND2_X1 i_34_80 (.A1(n_378), .A2(multiplicand[15]), .ZN(n_34_64));
   NAND4_X1 i_34_81 (.A1(n_34_61), .A2(n_34_62), .A3(n_34_63), .A4(n_34_64), 
      .ZN(n_395));
   NAND2_X1 i_34_82 (.A1(n_377), .A2(multiplicand[17]), .ZN(n_34_65));
   NAND2_X1 i_34_83 (.A1(n_375), .A2(n_64), .ZN(n_34_66));
   NAND2_X1 i_34_84 (.A1(n_376), .A2(n_63), .ZN(n_34_67));
   NAND2_X1 i_34_85 (.A1(n_378), .A2(multiplicand[16]), .ZN(n_34_68));
   NAND4_X1 i_34_86 (.A1(n_34_65), .A2(n_34_66), .A3(n_34_67), .A4(n_34_68), 
      .ZN(n_396));
   NAND2_X1 i_34_87 (.A1(n_377), .A2(multiplicand[18]), .ZN(n_34_69));
   NAND2_X1 i_34_88 (.A1(n_375), .A2(n_65), .ZN(n_34_70));
   NAND2_X1 i_34_89 (.A1(n_376), .A2(n_64), .ZN(n_34_71));
   NAND2_X1 i_34_90 (.A1(n_378), .A2(multiplicand[17]), .ZN(n_34_72));
   NAND4_X1 i_34_91 (.A1(n_34_69), .A2(n_34_70), .A3(n_34_71), .A4(n_34_72), 
      .ZN(n_397));
   NAND2_X1 i_34_92 (.A1(n_377), .A2(multiplicand[19]), .ZN(n_34_73));
   NAND2_X1 i_34_93 (.A1(n_375), .A2(n_66), .ZN(n_34_74));
   NAND2_X1 i_34_94 (.A1(n_376), .A2(n_65), .ZN(n_34_75));
   NAND2_X1 i_34_95 (.A1(n_378), .A2(multiplicand[18]), .ZN(n_34_76));
   NAND4_X1 i_34_96 (.A1(n_34_73), .A2(n_34_74), .A3(n_34_75), .A4(n_34_76), 
      .ZN(n_398));
   NAND2_X1 i_34_97 (.A1(n_377), .A2(multiplicand[20]), .ZN(n_34_77));
   NAND2_X1 i_34_98 (.A1(n_375), .A2(n_67), .ZN(n_34_78));
   NAND2_X1 i_34_99 (.A1(n_376), .A2(n_66), .ZN(n_34_79));
   NAND2_X1 i_34_100 (.A1(n_378), .A2(multiplicand[19]), .ZN(n_34_80));
   NAND4_X1 i_34_101 (.A1(n_34_77), .A2(n_34_78), .A3(n_34_79), .A4(n_34_80), 
      .ZN(n_399));
   NAND2_X1 i_34_102 (.A1(n_377), .A2(multiplicand[21]), .ZN(n_34_81));
   NAND2_X1 i_34_103 (.A1(n_375), .A2(n_68), .ZN(n_34_82));
   NAND2_X1 i_34_104 (.A1(n_376), .A2(n_67), .ZN(n_34_83));
   NAND2_X1 i_34_105 (.A1(n_378), .A2(multiplicand[20]), .ZN(n_34_84));
   NAND4_X1 i_34_106 (.A1(n_34_81), .A2(n_34_82), .A3(n_34_83), .A4(n_34_84), 
      .ZN(n_400));
   NAND2_X1 i_34_107 (.A1(n_377), .A2(multiplicand[22]), .ZN(n_34_85));
   NAND2_X1 i_34_108 (.A1(n_375), .A2(n_69), .ZN(n_34_86));
   NAND2_X1 i_34_109 (.A1(n_376), .A2(n_68), .ZN(n_34_87));
   NAND2_X1 i_34_110 (.A1(n_378), .A2(multiplicand[21]), .ZN(n_34_88));
   NAND4_X1 i_34_111 (.A1(n_34_85), .A2(n_34_86), .A3(n_34_87), .A4(n_34_88), 
      .ZN(n_401));
   NAND2_X1 i_34_112 (.A1(n_377), .A2(multiplicand[23]), .ZN(n_34_89));
   NAND2_X1 i_34_113 (.A1(n_375), .A2(n_70), .ZN(n_34_90));
   NAND2_X1 i_34_114 (.A1(n_376), .A2(n_69), .ZN(n_34_91));
   NAND2_X1 i_34_115 (.A1(n_378), .A2(multiplicand[22]), .ZN(n_34_92));
   NAND4_X1 i_34_116 (.A1(n_34_89), .A2(n_34_90), .A3(n_34_91), .A4(n_34_92), 
      .ZN(n_402));
   NAND2_X1 i_34_117 (.A1(n_377), .A2(multiplicand[24]), .ZN(n_34_93));
   NAND2_X1 i_34_118 (.A1(n_375), .A2(n_71), .ZN(n_34_94));
   NAND2_X1 i_34_119 (.A1(n_376), .A2(n_70), .ZN(n_34_95));
   NAND2_X1 i_34_120 (.A1(n_378), .A2(multiplicand[23]), .ZN(n_34_96));
   NAND4_X1 i_34_121 (.A1(n_34_93), .A2(n_34_94), .A3(n_34_95), .A4(n_34_96), 
      .ZN(n_403));
   NAND2_X1 i_34_122 (.A1(n_377), .A2(multiplicand[25]), .ZN(n_34_97));
   NAND2_X1 i_34_123 (.A1(n_375), .A2(n_72), .ZN(n_34_98));
   NAND2_X1 i_34_124 (.A1(n_376), .A2(n_71), .ZN(n_34_99));
   NAND2_X1 i_34_125 (.A1(n_378), .A2(multiplicand[24]), .ZN(n_34_100));
   NAND4_X1 i_34_126 (.A1(n_34_97), .A2(n_34_98), .A3(n_34_99), .A4(n_34_100), 
      .ZN(n_404));
   NAND2_X1 i_34_127 (.A1(n_377), .A2(multiplicand[26]), .ZN(n_34_101));
   NAND2_X1 i_34_128 (.A1(n_375), .A2(n_73), .ZN(n_34_102));
   NAND2_X1 i_34_129 (.A1(n_376), .A2(n_72), .ZN(n_34_103));
   NAND2_X1 i_34_130 (.A1(n_378), .A2(multiplicand[25]), .ZN(n_34_104));
   NAND4_X1 i_34_131 (.A1(n_34_101), .A2(n_34_102), .A3(n_34_103), .A4(n_34_104), 
      .ZN(n_405));
   NAND2_X1 i_34_132 (.A1(n_377), .A2(multiplicand[27]), .ZN(n_34_105));
   NAND2_X1 i_34_133 (.A1(n_375), .A2(n_74), .ZN(n_34_106));
   NAND2_X1 i_34_134 (.A1(n_376), .A2(n_73), .ZN(n_34_107));
   NAND2_X1 i_34_135 (.A1(n_378), .A2(multiplicand[26]), .ZN(n_34_108));
   NAND4_X1 i_34_136 (.A1(n_34_105), .A2(n_34_106), .A3(n_34_107), .A4(n_34_108), 
      .ZN(n_406));
   NAND2_X1 i_34_137 (.A1(n_377), .A2(multiplicand[28]), .ZN(n_34_109));
   NAND2_X1 i_34_138 (.A1(n_375), .A2(n_75), .ZN(n_34_110));
   NAND2_X1 i_34_139 (.A1(n_376), .A2(n_74), .ZN(n_34_111));
   NAND2_X1 i_34_140 (.A1(n_378), .A2(multiplicand[27]), .ZN(n_34_112));
   NAND4_X1 i_34_141 (.A1(n_34_109), .A2(n_34_110), .A3(n_34_111), .A4(n_34_112), 
      .ZN(n_407));
   NAND2_X1 i_34_142 (.A1(n_377), .A2(multiplicand[29]), .ZN(n_34_113));
   NAND2_X1 i_34_143 (.A1(n_375), .A2(n_76), .ZN(n_34_114));
   NAND2_X1 i_34_144 (.A1(n_376), .A2(n_75), .ZN(n_34_115));
   NAND2_X1 i_34_145 (.A1(n_378), .A2(multiplicand[28]), .ZN(n_34_116));
   NAND4_X1 i_34_146 (.A1(n_34_113), .A2(n_34_114), .A3(n_34_115), .A4(n_34_116), 
      .ZN(n_408));
   NAND2_X1 i_34_147 (.A1(n_377), .A2(multiplicand[30]), .ZN(n_34_117));
   NAND2_X1 i_34_148 (.A1(n_375), .A2(n_77), .ZN(n_34_118));
   NAND2_X1 i_34_149 (.A1(n_376), .A2(n_76), .ZN(n_34_119));
   NAND2_X1 i_34_150 (.A1(n_378), .A2(multiplicand[29]), .ZN(n_34_120));
   NAND4_X1 i_34_151 (.A1(n_34_117), .A2(n_34_118), .A3(n_34_119), .A4(n_34_120), 
      .ZN(n_409));
   NAND2_X1 i_34_152 (.A1(n_377), .A2(multiplicand[31]), .ZN(n_34_121));
   NAND2_X1 i_34_153 (.A1(n_375), .A2(n_78), .ZN(n_34_122));
   NAND2_X1 i_34_154 (.A1(n_376), .A2(n_77), .ZN(n_34_123));
   NAND2_X1 i_34_155 (.A1(n_378), .A2(multiplicand[30]), .ZN(n_34_124));
   NAND4_X1 i_34_156 (.A1(n_34_121), .A2(n_34_122), .A3(n_34_123), .A4(n_34_124), 
      .ZN(n_410));
   NAND2_X1 i_34_157 (.A1(n_376), .A2(n_78), .ZN(n_34_125));
   NAND2_X1 i_34_158 (.A1(n_378), .A2(multiplicand[31]), .ZN(n_34_126));
   NAND4_X1 i_34_159 (.A1(n_34_121), .A2(n_34_122), .A3(n_34_125), .A4(n_34_126), 
      .ZN(n_411));
   INV_X1 i_35_0 (.A(n_27), .ZN(n_35_0));
   AND3_X1 i_35_1 (.A1(n_35_0), .A2(n_28), .A3(n_29), .ZN(n_412));
   INV_X1 i_35_2 (.A(n_28), .ZN(n_35_1));
   AND3_X1 i_35_3 (.A1(n_35_1), .A2(n_27), .A3(n_29), .ZN(n_413));
   NOR3_X1 i_35_4 (.A1(n_35_1), .A2(n_27), .A3(n_29), .ZN(n_414));
   NOR3_X1 i_35_5 (.A1(n_35_0), .A2(n_28), .A3(n_29), .ZN(n_415));
   AOI22_X1 i_36_0 (.A1(n_414), .A2(multiplicand[0]), .B1(n_412), .B2(
      multiplicand[0]), .ZN(n_36_0));
   INV_X1 i_36_1 (.A(n_36_0), .ZN(n_416));
   NAND2_X1 i_36_2 (.A1(n_414), .A2(multiplicand[1]), .ZN(n_36_1));
   NAND2_X1 i_36_3 (.A1(n_412), .A2(n_48), .ZN(n_36_2));
   NAND2_X1 i_36_4 (.A1(n_413), .A2(multiplicand[0]), .ZN(n_36_3));
   NAND2_X1 i_36_5 (.A1(n_415), .A2(multiplicand[0]), .ZN(n_36_4));
   NAND4_X1 i_36_6 (.A1(n_36_1), .A2(n_36_2), .A3(n_36_3), .A4(n_36_4), .ZN(
      n_417));
   NAND2_X1 i_36_7 (.A1(n_414), .A2(multiplicand[2]), .ZN(n_36_5));
   NAND2_X1 i_36_8 (.A1(n_412), .A2(n_49), .ZN(n_36_6));
   NAND2_X1 i_36_9 (.A1(n_413), .A2(n_48), .ZN(n_36_7));
   NAND2_X1 i_36_10 (.A1(n_415), .A2(multiplicand[1]), .ZN(n_36_8));
   NAND4_X1 i_36_11 (.A1(n_36_5), .A2(n_36_6), .A3(n_36_7), .A4(n_36_8), 
      .ZN(n_418));
   NAND2_X1 i_36_12 (.A1(n_414), .A2(multiplicand[3]), .ZN(n_36_9));
   NAND2_X1 i_36_13 (.A1(n_412), .A2(n_50), .ZN(n_36_10));
   NAND2_X1 i_36_14 (.A1(n_413), .A2(n_49), .ZN(n_36_11));
   NAND2_X1 i_36_15 (.A1(n_415), .A2(multiplicand[2]), .ZN(n_36_12));
   NAND4_X1 i_36_16 (.A1(n_36_9), .A2(n_36_10), .A3(n_36_11), .A4(n_36_12), 
      .ZN(n_419));
   NAND2_X1 i_36_17 (.A1(n_414), .A2(multiplicand[4]), .ZN(n_36_13));
   NAND2_X1 i_36_18 (.A1(n_412), .A2(n_51), .ZN(n_36_14));
   NAND2_X1 i_36_19 (.A1(n_413), .A2(n_50), .ZN(n_36_15));
   NAND2_X1 i_36_20 (.A1(n_415), .A2(multiplicand[3]), .ZN(n_36_16));
   NAND4_X1 i_36_21 (.A1(n_36_13), .A2(n_36_14), .A3(n_36_15), .A4(n_36_16), 
      .ZN(n_420));
   NAND2_X1 i_36_22 (.A1(n_414), .A2(multiplicand[5]), .ZN(n_36_17));
   NAND2_X1 i_36_23 (.A1(n_412), .A2(n_52), .ZN(n_36_18));
   NAND2_X1 i_36_24 (.A1(n_413), .A2(n_51), .ZN(n_36_19));
   NAND2_X1 i_36_25 (.A1(n_415), .A2(multiplicand[4]), .ZN(n_36_20));
   NAND4_X1 i_36_26 (.A1(n_36_17), .A2(n_36_18), .A3(n_36_19), .A4(n_36_20), 
      .ZN(n_421));
   NAND2_X1 i_36_27 (.A1(n_414), .A2(multiplicand[6]), .ZN(n_36_21));
   NAND2_X1 i_36_28 (.A1(n_412), .A2(n_53), .ZN(n_36_22));
   NAND2_X1 i_36_29 (.A1(n_413), .A2(n_52), .ZN(n_36_23));
   NAND2_X1 i_36_30 (.A1(n_415), .A2(multiplicand[5]), .ZN(n_36_24));
   NAND4_X1 i_36_31 (.A1(n_36_21), .A2(n_36_22), .A3(n_36_23), .A4(n_36_24), 
      .ZN(n_422));
   NAND2_X1 i_36_32 (.A1(n_414), .A2(multiplicand[7]), .ZN(n_36_25));
   NAND2_X1 i_36_33 (.A1(n_412), .A2(n_54), .ZN(n_36_26));
   NAND2_X1 i_36_34 (.A1(n_413), .A2(n_53), .ZN(n_36_27));
   NAND2_X1 i_36_35 (.A1(n_415), .A2(multiplicand[6]), .ZN(n_36_28));
   NAND4_X1 i_36_36 (.A1(n_36_25), .A2(n_36_26), .A3(n_36_27), .A4(n_36_28), 
      .ZN(n_423));
   NAND2_X1 i_36_37 (.A1(n_414), .A2(multiplicand[8]), .ZN(n_36_29));
   NAND2_X1 i_36_38 (.A1(n_412), .A2(n_55), .ZN(n_36_30));
   NAND2_X1 i_36_39 (.A1(n_413), .A2(n_54), .ZN(n_36_31));
   NAND2_X1 i_36_40 (.A1(n_415), .A2(multiplicand[7]), .ZN(n_36_32));
   NAND4_X1 i_36_41 (.A1(n_36_29), .A2(n_36_30), .A3(n_36_31), .A4(n_36_32), 
      .ZN(n_424));
   NAND2_X1 i_36_42 (.A1(n_414), .A2(multiplicand[9]), .ZN(n_36_33));
   NAND2_X1 i_36_43 (.A1(n_412), .A2(n_56), .ZN(n_36_34));
   NAND2_X1 i_36_44 (.A1(n_413), .A2(n_55), .ZN(n_36_35));
   NAND2_X1 i_36_45 (.A1(n_415), .A2(multiplicand[8]), .ZN(n_36_36));
   NAND4_X1 i_36_46 (.A1(n_36_33), .A2(n_36_34), .A3(n_36_35), .A4(n_36_36), 
      .ZN(n_425));
   NAND2_X1 i_36_47 (.A1(n_414), .A2(multiplicand[10]), .ZN(n_36_37));
   NAND2_X1 i_36_48 (.A1(n_412), .A2(n_57), .ZN(n_36_38));
   NAND2_X1 i_36_49 (.A1(n_413), .A2(n_56), .ZN(n_36_39));
   NAND2_X1 i_36_50 (.A1(n_415), .A2(multiplicand[9]), .ZN(n_36_40));
   NAND4_X1 i_36_51 (.A1(n_36_37), .A2(n_36_38), .A3(n_36_39), .A4(n_36_40), 
      .ZN(n_426));
   NAND2_X1 i_36_52 (.A1(n_414), .A2(multiplicand[11]), .ZN(n_36_41));
   NAND2_X1 i_36_53 (.A1(n_412), .A2(n_58), .ZN(n_36_42));
   NAND2_X1 i_36_54 (.A1(n_413), .A2(n_57), .ZN(n_36_43));
   NAND2_X1 i_36_55 (.A1(n_415), .A2(multiplicand[10]), .ZN(n_36_44));
   NAND4_X1 i_36_56 (.A1(n_36_41), .A2(n_36_42), .A3(n_36_43), .A4(n_36_44), 
      .ZN(n_427));
   NAND2_X1 i_36_57 (.A1(n_414), .A2(multiplicand[12]), .ZN(n_36_45));
   NAND2_X1 i_36_58 (.A1(n_412), .A2(n_59), .ZN(n_36_46));
   NAND2_X1 i_36_59 (.A1(n_413), .A2(n_58), .ZN(n_36_47));
   NAND2_X1 i_36_60 (.A1(n_415), .A2(multiplicand[11]), .ZN(n_36_48));
   NAND4_X1 i_36_61 (.A1(n_36_45), .A2(n_36_46), .A3(n_36_47), .A4(n_36_48), 
      .ZN(n_428));
   NAND2_X1 i_36_62 (.A1(n_414), .A2(multiplicand[13]), .ZN(n_36_49));
   NAND2_X1 i_36_63 (.A1(n_412), .A2(n_60), .ZN(n_36_50));
   NAND2_X1 i_36_64 (.A1(n_413), .A2(n_59), .ZN(n_36_51));
   NAND2_X1 i_36_65 (.A1(n_415), .A2(multiplicand[12]), .ZN(n_36_52));
   NAND4_X1 i_36_66 (.A1(n_36_49), .A2(n_36_50), .A3(n_36_51), .A4(n_36_52), 
      .ZN(n_429));
   NAND2_X1 i_36_67 (.A1(n_414), .A2(multiplicand[14]), .ZN(n_36_53));
   NAND2_X1 i_36_68 (.A1(n_412), .A2(n_61), .ZN(n_36_54));
   NAND2_X1 i_36_69 (.A1(n_413), .A2(n_60), .ZN(n_36_55));
   NAND2_X1 i_36_70 (.A1(n_415), .A2(multiplicand[13]), .ZN(n_36_56));
   NAND4_X1 i_36_71 (.A1(n_36_53), .A2(n_36_54), .A3(n_36_55), .A4(n_36_56), 
      .ZN(n_430));
   NAND2_X1 i_36_72 (.A1(n_414), .A2(multiplicand[15]), .ZN(n_36_57));
   NAND2_X1 i_36_73 (.A1(n_412), .A2(n_62), .ZN(n_36_58));
   NAND2_X1 i_36_74 (.A1(n_413), .A2(n_61), .ZN(n_36_59));
   NAND2_X1 i_36_75 (.A1(n_415), .A2(multiplicand[14]), .ZN(n_36_60));
   NAND4_X1 i_36_76 (.A1(n_36_57), .A2(n_36_58), .A3(n_36_59), .A4(n_36_60), 
      .ZN(n_431));
   NAND2_X1 i_36_77 (.A1(n_414), .A2(multiplicand[16]), .ZN(n_36_61));
   NAND2_X1 i_36_78 (.A1(n_412), .A2(n_63), .ZN(n_36_62));
   NAND2_X1 i_36_79 (.A1(n_413), .A2(n_62), .ZN(n_36_63));
   NAND2_X1 i_36_80 (.A1(n_415), .A2(multiplicand[15]), .ZN(n_36_64));
   NAND4_X1 i_36_81 (.A1(n_36_61), .A2(n_36_62), .A3(n_36_63), .A4(n_36_64), 
      .ZN(n_432));
   NAND2_X1 i_36_82 (.A1(n_414), .A2(multiplicand[17]), .ZN(n_36_65));
   NAND2_X1 i_36_83 (.A1(n_412), .A2(n_64), .ZN(n_36_66));
   NAND2_X1 i_36_84 (.A1(n_413), .A2(n_63), .ZN(n_36_67));
   NAND2_X1 i_36_85 (.A1(n_415), .A2(multiplicand[16]), .ZN(n_36_68));
   NAND4_X1 i_36_86 (.A1(n_36_65), .A2(n_36_66), .A3(n_36_67), .A4(n_36_68), 
      .ZN(n_433));
   NAND2_X1 i_36_87 (.A1(n_414), .A2(multiplicand[18]), .ZN(n_36_69));
   NAND2_X1 i_36_88 (.A1(n_412), .A2(n_65), .ZN(n_36_70));
   NAND2_X1 i_36_89 (.A1(n_413), .A2(n_64), .ZN(n_36_71));
   NAND2_X1 i_36_90 (.A1(n_415), .A2(multiplicand[17]), .ZN(n_36_72));
   NAND4_X1 i_36_91 (.A1(n_36_69), .A2(n_36_70), .A3(n_36_71), .A4(n_36_72), 
      .ZN(n_434));
   NAND2_X1 i_36_92 (.A1(n_414), .A2(multiplicand[19]), .ZN(n_36_73));
   NAND2_X1 i_36_93 (.A1(n_412), .A2(n_66), .ZN(n_36_74));
   NAND2_X1 i_36_94 (.A1(n_413), .A2(n_65), .ZN(n_36_75));
   NAND2_X1 i_36_95 (.A1(n_415), .A2(multiplicand[18]), .ZN(n_36_76));
   NAND4_X1 i_36_96 (.A1(n_36_73), .A2(n_36_74), .A3(n_36_75), .A4(n_36_76), 
      .ZN(n_435));
   NAND2_X1 i_36_97 (.A1(n_414), .A2(multiplicand[20]), .ZN(n_36_77));
   NAND2_X1 i_36_98 (.A1(n_412), .A2(n_67), .ZN(n_36_78));
   NAND2_X1 i_36_99 (.A1(n_413), .A2(n_66), .ZN(n_36_79));
   NAND2_X1 i_36_100 (.A1(n_415), .A2(multiplicand[19]), .ZN(n_36_80));
   NAND4_X1 i_36_101 (.A1(n_36_77), .A2(n_36_78), .A3(n_36_79), .A4(n_36_80), 
      .ZN(n_436));
   NAND2_X1 i_36_102 (.A1(n_414), .A2(multiplicand[21]), .ZN(n_36_81));
   NAND2_X1 i_36_103 (.A1(n_412), .A2(n_68), .ZN(n_36_82));
   NAND2_X1 i_36_104 (.A1(n_413), .A2(n_67), .ZN(n_36_83));
   NAND2_X1 i_36_105 (.A1(n_415), .A2(multiplicand[20]), .ZN(n_36_84));
   NAND4_X1 i_36_106 (.A1(n_36_81), .A2(n_36_82), .A3(n_36_83), .A4(n_36_84), 
      .ZN(n_437));
   NAND2_X1 i_36_107 (.A1(n_414), .A2(multiplicand[22]), .ZN(n_36_85));
   NAND2_X1 i_36_108 (.A1(n_412), .A2(n_69), .ZN(n_36_86));
   NAND2_X1 i_36_109 (.A1(n_413), .A2(n_68), .ZN(n_36_87));
   NAND2_X1 i_36_110 (.A1(n_415), .A2(multiplicand[21]), .ZN(n_36_88));
   NAND4_X1 i_36_111 (.A1(n_36_85), .A2(n_36_86), .A3(n_36_87), .A4(n_36_88), 
      .ZN(n_438));
   NAND2_X1 i_36_112 (.A1(n_414), .A2(multiplicand[23]), .ZN(n_36_89));
   NAND2_X1 i_36_113 (.A1(n_412), .A2(n_70), .ZN(n_36_90));
   NAND2_X1 i_36_114 (.A1(n_413), .A2(n_69), .ZN(n_36_91));
   NAND2_X1 i_36_115 (.A1(n_415), .A2(multiplicand[22]), .ZN(n_36_92));
   NAND4_X1 i_36_116 (.A1(n_36_89), .A2(n_36_90), .A3(n_36_91), .A4(n_36_92), 
      .ZN(n_439));
   NAND2_X1 i_36_117 (.A1(n_414), .A2(multiplicand[24]), .ZN(n_36_93));
   NAND2_X1 i_36_118 (.A1(n_412), .A2(n_71), .ZN(n_36_94));
   NAND2_X1 i_36_119 (.A1(n_413), .A2(n_70), .ZN(n_36_95));
   NAND2_X1 i_36_120 (.A1(n_415), .A2(multiplicand[23]), .ZN(n_36_96));
   NAND4_X1 i_36_121 (.A1(n_36_93), .A2(n_36_94), .A3(n_36_95), .A4(n_36_96), 
      .ZN(n_440));
   NAND2_X1 i_36_122 (.A1(n_414), .A2(multiplicand[25]), .ZN(n_36_97));
   NAND2_X1 i_36_123 (.A1(n_412), .A2(n_72), .ZN(n_36_98));
   NAND2_X1 i_36_124 (.A1(n_413), .A2(n_71), .ZN(n_36_99));
   NAND2_X1 i_36_125 (.A1(n_415), .A2(multiplicand[24]), .ZN(n_36_100));
   NAND4_X1 i_36_126 (.A1(n_36_97), .A2(n_36_98), .A3(n_36_99), .A4(n_36_100), 
      .ZN(n_441));
   NAND2_X1 i_36_127 (.A1(n_414), .A2(multiplicand[26]), .ZN(n_36_101));
   NAND2_X1 i_36_128 (.A1(n_412), .A2(n_73), .ZN(n_36_102));
   NAND2_X1 i_36_129 (.A1(n_413), .A2(n_72), .ZN(n_36_103));
   NAND2_X1 i_36_130 (.A1(n_415), .A2(multiplicand[25]), .ZN(n_36_104));
   NAND4_X1 i_36_131 (.A1(n_36_101), .A2(n_36_102), .A3(n_36_103), .A4(n_36_104), 
      .ZN(n_442));
   NAND2_X1 i_36_132 (.A1(n_414), .A2(multiplicand[27]), .ZN(n_36_105));
   NAND2_X1 i_36_133 (.A1(n_412), .A2(n_74), .ZN(n_36_106));
   NAND2_X1 i_36_134 (.A1(n_413), .A2(n_73), .ZN(n_36_107));
   NAND2_X1 i_36_135 (.A1(n_415), .A2(multiplicand[26]), .ZN(n_36_108));
   NAND4_X1 i_36_136 (.A1(n_36_105), .A2(n_36_106), .A3(n_36_107), .A4(n_36_108), 
      .ZN(n_443));
   NAND2_X1 i_36_137 (.A1(n_414), .A2(multiplicand[28]), .ZN(n_36_109));
   NAND2_X1 i_36_138 (.A1(n_412), .A2(n_75), .ZN(n_36_110));
   NAND2_X1 i_36_139 (.A1(n_413), .A2(n_74), .ZN(n_36_111));
   NAND2_X1 i_36_140 (.A1(n_415), .A2(multiplicand[27]), .ZN(n_36_112));
   NAND4_X1 i_36_141 (.A1(n_36_109), .A2(n_36_110), .A3(n_36_111), .A4(n_36_112), 
      .ZN(n_444));
   NAND2_X1 i_36_142 (.A1(n_414), .A2(multiplicand[29]), .ZN(n_36_113));
   NAND2_X1 i_36_143 (.A1(n_412), .A2(n_76), .ZN(n_36_114));
   NAND2_X1 i_36_144 (.A1(n_413), .A2(n_75), .ZN(n_36_115));
   NAND2_X1 i_36_145 (.A1(n_415), .A2(multiplicand[28]), .ZN(n_36_116));
   NAND4_X1 i_36_146 (.A1(n_36_113), .A2(n_36_114), .A3(n_36_115), .A4(n_36_116), 
      .ZN(n_445));
   NAND2_X1 i_36_147 (.A1(n_414), .A2(multiplicand[30]), .ZN(n_36_117));
   NAND2_X1 i_36_148 (.A1(n_412), .A2(n_77), .ZN(n_36_118));
   NAND2_X1 i_36_149 (.A1(n_413), .A2(n_76), .ZN(n_36_119));
   NAND2_X1 i_36_150 (.A1(n_415), .A2(multiplicand[29]), .ZN(n_36_120));
   NAND4_X1 i_36_151 (.A1(n_36_117), .A2(n_36_118), .A3(n_36_119), .A4(n_36_120), 
      .ZN(n_446));
   NAND2_X1 i_36_152 (.A1(n_414), .A2(multiplicand[31]), .ZN(n_36_121));
   NAND2_X1 i_36_153 (.A1(n_412), .A2(n_78), .ZN(n_36_122));
   NAND2_X1 i_36_154 (.A1(n_413), .A2(n_77), .ZN(n_36_123));
   NAND2_X1 i_36_155 (.A1(n_415), .A2(multiplicand[30]), .ZN(n_36_124));
   NAND4_X1 i_36_156 (.A1(n_36_121), .A2(n_36_122), .A3(n_36_123), .A4(n_36_124), 
      .ZN(n_447));
   NAND2_X1 i_36_157 (.A1(n_413), .A2(n_78), .ZN(n_36_125));
   NAND2_X1 i_36_158 (.A1(n_415), .A2(multiplicand[31]), .ZN(n_36_126));
   NAND4_X1 i_36_159 (.A1(n_36_121), .A2(n_36_122), .A3(n_36_125), .A4(n_36_126), 
      .ZN(n_448));
   INV_X1 i_37_0 (.A(n_30), .ZN(n_37_0));
   AND3_X1 i_37_1 (.A1(n_37_0), .A2(n_31), .A3(n_32), .ZN(n_449));
   INV_X1 i_37_2 (.A(n_31), .ZN(n_37_1));
   AND3_X1 i_37_3 (.A1(n_37_1), .A2(n_30), .A3(n_32), .ZN(n_450));
   NOR3_X1 i_37_4 (.A1(n_37_1), .A2(n_30), .A3(n_32), .ZN(n_451));
   NOR3_X1 i_37_5 (.A1(n_37_0), .A2(n_31), .A3(n_32), .ZN(n_452));
   AOI22_X1 i_38_0 (.A1(n_451), .A2(multiplicand[0]), .B1(n_449), .B2(
      multiplicand[0]), .ZN(n_38_0));
   INV_X1 i_38_1 (.A(n_38_0), .ZN(n_453));
   NAND2_X1 i_38_2 (.A1(n_451), .A2(multiplicand[1]), .ZN(n_38_1));
   NAND2_X1 i_38_3 (.A1(n_449), .A2(n_48), .ZN(n_38_2));
   NAND2_X1 i_38_4 (.A1(n_450), .A2(multiplicand[0]), .ZN(n_38_3));
   NAND2_X1 i_38_5 (.A1(n_452), .A2(multiplicand[0]), .ZN(n_38_4));
   NAND4_X1 i_38_6 (.A1(n_38_1), .A2(n_38_2), .A3(n_38_3), .A4(n_38_4), .ZN(
      n_454));
   NAND2_X1 i_38_7 (.A1(n_451), .A2(multiplicand[2]), .ZN(n_38_5));
   NAND2_X1 i_38_8 (.A1(n_449), .A2(n_49), .ZN(n_38_6));
   NAND2_X1 i_38_9 (.A1(n_450), .A2(n_48), .ZN(n_38_7));
   NAND2_X1 i_38_10 (.A1(n_452), .A2(multiplicand[1]), .ZN(n_38_8));
   NAND4_X1 i_38_11 (.A1(n_38_5), .A2(n_38_6), .A3(n_38_7), .A4(n_38_8), 
      .ZN(n_455));
   NAND2_X1 i_38_12 (.A1(n_451), .A2(multiplicand[3]), .ZN(n_38_9));
   NAND2_X1 i_38_13 (.A1(n_449), .A2(n_50), .ZN(n_38_10));
   NAND2_X1 i_38_14 (.A1(n_450), .A2(n_49), .ZN(n_38_11));
   NAND2_X1 i_38_15 (.A1(n_452), .A2(multiplicand[2]), .ZN(n_38_12));
   NAND4_X1 i_38_16 (.A1(n_38_9), .A2(n_38_10), .A3(n_38_11), .A4(n_38_12), 
      .ZN(n_456));
   NAND2_X1 i_38_17 (.A1(n_451), .A2(multiplicand[4]), .ZN(n_38_13));
   NAND2_X1 i_38_18 (.A1(n_449), .A2(n_51), .ZN(n_38_14));
   NAND2_X1 i_38_19 (.A1(n_450), .A2(n_50), .ZN(n_38_15));
   NAND2_X1 i_38_20 (.A1(n_452), .A2(multiplicand[3]), .ZN(n_38_16));
   NAND4_X1 i_38_21 (.A1(n_38_13), .A2(n_38_14), .A3(n_38_15), .A4(n_38_16), 
      .ZN(n_457));
   NAND2_X1 i_38_22 (.A1(n_451), .A2(multiplicand[5]), .ZN(n_38_17));
   NAND2_X1 i_38_23 (.A1(n_449), .A2(n_52), .ZN(n_38_18));
   NAND2_X1 i_38_24 (.A1(n_450), .A2(n_51), .ZN(n_38_19));
   NAND2_X1 i_38_25 (.A1(n_452), .A2(multiplicand[4]), .ZN(n_38_20));
   NAND4_X1 i_38_26 (.A1(n_38_17), .A2(n_38_18), .A3(n_38_19), .A4(n_38_20), 
      .ZN(n_458));
   NAND2_X1 i_38_27 (.A1(n_451), .A2(multiplicand[6]), .ZN(n_38_21));
   NAND2_X1 i_38_28 (.A1(n_449), .A2(n_53), .ZN(n_38_22));
   NAND2_X1 i_38_29 (.A1(n_450), .A2(n_52), .ZN(n_38_23));
   NAND2_X1 i_38_30 (.A1(n_452), .A2(multiplicand[5]), .ZN(n_38_24));
   NAND4_X1 i_38_31 (.A1(n_38_21), .A2(n_38_22), .A3(n_38_23), .A4(n_38_24), 
      .ZN(n_459));
   NAND2_X1 i_38_32 (.A1(n_451), .A2(multiplicand[7]), .ZN(n_38_25));
   NAND2_X1 i_38_33 (.A1(n_449), .A2(n_54), .ZN(n_38_26));
   NAND2_X1 i_38_34 (.A1(n_450), .A2(n_53), .ZN(n_38_27));
   NAND2_X1 i_38_35 (.A1(n_452), .A2(multiplicand[6]), .ZN(n_38_28));
   NAND4_X1 i_38_36 (.A1(n_38_25), .A2(n_38_26), .A3(n_38_27), .A4(n_38_28), 
      .ZN(n_460));
   NAND2_X1 i_38_37 (.A1(n_451), .A2(multiplicand[8]), .ZN(n_38_29));
   NAND2_X1 i_38_38 (.A1(n_449), .A2(n_55), .ZN(n_38_30));
   NAND2_X1 i_38_39 (.A1(n_450), .A2(n_54), .ZN(n_38_31));
   NAND2_X1 i_38_40 (.A1(n_452), .A2(multiplicand[7]), .ZN(n_38_32));
   NAND4_X1 i_38_41 (.A1(n_38_29), .A2(n_38_30), .A3(n_38_31), .A4(n_38_32), 
      .ZN(n_461));
   NAND2_X1 i_38_42 (.A1(n_451), .A2(multiplicand[9]), .ZN(n_38_33));
   NAND2_X1 i_38_43 (.A1(n_449), .A2(n_56), .ZN(n_38_34));
   NAND2_X1 i_38_44 (.A1(n_450), .A2(n_55), .ZN(n_38_35));
   NAND2_X1 i_38_45 (.A1(n_452), .A2(multiplicand[8]), .ZN(n_38_36));
   NAND4_X1 i_38_46 (.A1(n_38_33), .A2(n_38_34), .A3(n_38_35), .A4(n_38_36), 
      .ZN(n_462));
   NAND2_X1 i_38_47 (.A1(n_451), .A2(multiplicand[10]), .ZN(n_38_37));
   NAND2_X1 i_38_48 (.A1(n_449), .A2(n_57), .ZN(n_38_38));
   NAND2_X1 i_38_49 (.A1(n_450), .A2(n_56), .ZN(n_38_39));
   NAND2_X1 i_38_50 (.A1(n_452), .A2(multiplicand[9]), .ZN(n_38_40));
   NAND4_X1 i_38_51 (.A1(n_38_37), .A2(n_38_38), .A3(n_38_39), .A4(n_38_40), 
      .ZN(n_463));
   NAND2_X1 i_38_52 (.A1(n_451), .A2(multiplicand[11]), .ZN(n_38_41));
   NAND2_X1 i_38_53 (.A1(n_449), .A2(n_58), .ZN(n_38_42));
   NAND2_X1 i_38_54 (.A1(n_450), .A2(n_57), .ZN(n_38_43));
   NAND2_X1 i_38_55 (.A1(n_452), .A2(multiplicand[10]), .ZN(n_38_44));
   NAND4_X1 i_38_56 (.A1(n_38_41), .A2(n_38_42), .A3(n_38_43), .A4(n_38_44), 
      .ZN(n_464));
   NAND2_X1 i_38_57 (.A1(n_451), .A2(multiplicand[12]), .ZN(n_38_45));
   NAND2_X1 i_38_58 (.A1(n_449), .A2(n_59), .ZN(n_38_46));
   NAND2_X1 i_38_59 (.A1(n_450), .A2(n_58), .ZN(n_38_47));
   NAND2_X1 i_38_60 (.A1(n_452), .A2(multiplicand[11]), .ZN(n_38_48));
   NAND4_X1 i_38_61 (.A1(n_38_45), .A2(n_38_46), .A3(n_38_47), .A4(n_38_48), 
      .ZN(n_465));
   NAND2_X1 i_38_62 (.A1(n_451), .A2(multiplicand[13]), .ZN(n_38_49));
   NAND2_X1 i_38_63 (.A1(n_449), .A2(n_60), .ZN(n_38_50));
   NAND2_X1 i_38_64 (.A1(n_450), .A2(n_59), .ZN(n_38_51));
   NAND2_X1 i_38_65 (.A1(n_452), .A2(multiplicand[12]), .ZN(n_38_52));
   NAND4_X1 i_38_66 (.A1(n_38_49), .A2(n_38_50), .A3(n_38_51), .A4(n_38_52), 
      .ZN(n_466));
   NAND2_X1 i_38_67 (.A1(n_451), .A2(multiplicand[14]), .ZN(n_38_53));
   NAND2_X1 i_38_68 (.A1(n_449), .A2(n_61), .ZN(n_38_54));
   NAND2_X1 i_38_69 (.A1(n_450), .A2(n_60), .ZN(n_38_55));
   NAND2_X1 i_38_70 (.A1(n_452), .A2(multiplicand[13]), .ZN(n_38_56));
   NAND4_X1 i_38_71 (.A1(n_38_53), .A2(n_38_54), .A3(n_38_55), .A4(n_38_56), 
      .ZN(n_467));
   NAND2_X1 i_38_72 (.A1(n_451), .A2(multiplicand[15]), .ZN(n_38_57));
   NAND2_X1 i_38_73 (.A1(n_449), .A2(n_62), .ZN(n_38_58));
   NAND2_X1 i_38_74 (.A1(n_450), .A2(n_61), .ZN(n_38_59));
   NAND2_X1 i_38_75 (.A1(n_452), .A2(multiplicand[14]), .ZN(n_38_60));
   NAND4_X1 i_38_76 (.A1(n_38_57), .A2(n_38_58), .A3(n_38_59), .A4(n_38_60), 
      .ZN(n_468));
   NAND2_X1 i_38_77 (.A1(n_451), .A2(multiplicand[16]), .ZN(n_38_61));
   NAND2_X1 i_38_78 (.A1(n_449), .A2(n_63), .ZN(n_38_62));
   NAND2_X1 i_38_79 (.A1(n_450), .A2(n_62), .ZN(n_38_63));
   NAND2_X1 i_38_80 (.A1(n_452), .A2(multiplicand[15]), .ZN(n_38_64));
   NAND4_X1 i_38_81 (.A1(n_38_61), .A2(n_38_62), .A3(n_38_63), .A4(n_38_64), 
      .ZN(n_469));
   NAND2_X1 i_38_82 (.A1(n_451), .A2(multiplicand[17]), .ZN(n_38_65));
   NAND2_X1 i_38_83 (.A1(n_449), .A2(n_64), .ZN(n_38_66));
   NAND2_X1 i_38_84 (.A1(n_450), .A2(n_63), .ZN(n_38_67));
   NAND2_X1 i_38_85 (.A1(n_452), .A2(multiplicand[16]), .ZN(n_38_68));
   NAND4_X1 i_38_86 (.A1(n_38_65), .A2(n_38_66), .A3(n_38_67), .A4(n_38_68), 
      .ZN(n_470));
   NAND2_X1 i_38_87 (.A1(n_451), .A2(multiplicand[18]), .ZN(n_38_69));
   NAND2_X1 i_38_88 (.A1(n_449), .A2(n_65), .ZN(n_38_70));
   NAND2_X1 i_38_89 (.A1(n_450), .A2(n_64), .ZN(n_38_71));
   NAND2_X1 i_38_90 (.A1(n_452), .A2(multiplicand[17]), .ZN(n_38_72));
   NAND4_X1 i_38_91 (.A1(n_38_69), .A2(n_38_70), .A3(n_38_71), .A4(n_38_72), 
      .ZN(n_471));
   NAND2_X1 i_38_92 (.A1(n_451), .A2(multiplicand[19]), .ZN(n_38_73));
   NAND2_X1 i_38_93 (.A1(n_449), .A2(n_66), .ZN(n_38_74));
   NAND2_X1 i_38_94 (.A1(n_450), .A2(n_65), .ZN(n_38_75));
   NAND2_X1 i_38_95 (.A1(n_452), .A2(multiplicand[18]), .ZN(n_38_76));
   NAND4_X1 i_38_96 (.A1(n_38_73), .A2(n_38_74), .A3(n_38_75), .A4(n_38_76), 
      .ZN(n_472));
   NAND2_X1 i_38_97 (.A1(n_451), .A2(multiplicand[20]), .ZN(n_38_77));
   NAND2_X1 i_38_98 (.A1(n_449), .A2(n_67), .ZN(n_38_78));
   NAND2_X1 i_38_99 (.A1(n_450), .A2(n_66), .ZN(n_38_79));
   NAND2_X1 i_38_100 (.A1(n_452), .A2(multiplicand[19]), .ZN(n_38_80));
   NAND4_X1 i_38_101 (.A1(n_38_77), .A2(n_38_78), .A3(n_38_79), .A4(n_38_80), 
      .ZN(n_473));
   NAND2_X1 i_38_102 (.A1(n_451), .A2(multiplicand[21]), .ZN(n_38_81));
   NAND2_X1 i_38_103 (.A1(n_449), .A2(n_68), .ZN(n_38_82));
   NAND2_X1 i_38_104 (.A1(n_450), .A2(n_67), .ZN(n_38_83));
   NAND2_X1 i_38_105 (.A1(n_452), .A2(multiplicand[20]), .ZN(n_38_84));
   NAND4_X1 i_38_106 (.A1(n_38_81), .A2(n_38_82), .A3(n_38_83), .A4(n_38_84), 
      .ZN(n_474));
   NAND2_X1 i_38_107 (.A1(n_451), .A2(multiplicand[22]), .ZN(n_38_85));
   NAND2_X1 i_38_108 (.A1(n_449), .A2(n_69), .ZN(n_38_86));
   NAND2_X1 i_38_109 (.A1(n_450), .A2(n_68), .ZN(n_38_87));
   NAND2_X1 i_38_110 (.A1(n_452), .A2(multiplicand[21]), .ZN(n_38_88));
   NAND4_X1 i_38_111 (.A1(n_38_85), .A2(n_38_86), .A3(n_38_87), .A4(n_38_88), 
      .ZN(n_475));
   NAND2_X1 i_38_112 (.A1(n_451), .A2(multiplicand[23]), .ZN(n_38_89));
   NAND2_X1 i_38_113 (.A1(n_449), .A2(n_70), .ZN(n_38_90));
   NAND2_X1 i_38_114 (.A1(n_450), .A2(n_69), .ZN(n_38_91));
   NAND2_X1 i_38_115 (.A1(n_452), .A2(multiplicand[22]), .ZN(n_38_92));
   NAND4_X1 i_38_116 (.A1(n_38_89), .A2(n_38_90), .A3(n_38_91), .A4(n_38_92), 
      .ZN(n_476));
   NAND2_X1 i_38_117 (.A1(n_451), .A2(multiplicand[24]), .ZN(n_38_93));
   NAND2_X1 i_38_118 (.A1(n_449), .A2(n_71), .ZN(n_38_94));
   NAND2_X1 i_38_119 (.A1(n_450), .A2(n_70), .ZN(n_38_95));
   NAND2_X1 i_38_120 (.A1(n_452), .A2(multiplicand[23]), .ZN(n_38_96));
   NAND4_X1 i_38_121 (.A1(n_38_93), .A2(n_38_94), .A3(n_38_95), .A4(n_38_96), 
      .ZN(n_477));
   NAND2_X1 i_38_122 (.A1(n_451), .A2(multiplicand[25]), .ZN(n_38_97));
   NAND2_X1 i_38_123 (.A1(n_449), .A2(n_72), .ZN(n_38_98));
   NAND2_X1 i_38_124 (.A1(n_450), .A2(n_71), .ZN(n_38_99));
   NAND2_X1 i_38_125 (.A1(n_452), .A2(multiplicand[24]), .ZN(n_38_100));
   NAND4_X1 i_38_126 (.A1(n_38_97), .A2(n_38_98), .A3(n_38_99), .A4(n_38_100), 
      .ZN(n_478));
   NAND2_X1 i_38_127 (.A1(n_451), .A2(multiplicand[26]), .ZN(n_38_101));
   NAND2_X1 i_38_128 (.A1(n_449), .A2(n_73), .ZN(n_38_102));
   NAND2_X1 i_38_129 (.A1(n_450), .A2(n_72), .ZN(n_38_103));
   NAND2_X1 i_38_130 (.A1(n_452), .A2(multiplicand[25]), .ZN(n_38_104));
   NAND4_X1 i_38_131 (.A1(n_38_101), .A2(n_38_102), .A3(n_38_103), .A4(n_38_104), 
      .ZN(n_479));
   NAND2_X1 i_38_132 (.A1(n_451), .A2(multiplicand[27]), .ZN(n_38_105));
   NAND2_X1 i_38_133 (.A1(n_449), .A2(n_74), .ZN(n_38_106));
   NAND2_X1 i_38_134 (.A1(n_450), .A2(n_73), .ZN(n_38_107));
   NAND2_X1 i_38_135 (.A1(n_452), .A2(multiplicand[26]), .ZN(n_38_108));
   NAND4_X1 i_38_136 (.A1(n_38_105), .A2(n_38_106), .A3(n_38_107), .A4(n_38_108), 
      .ZN(n_480));
   NAND2_X1 i_38_137 (.A1(n_451), .A2(multiplicand[28]), .ZN(n_38_109));
   NAND2_X1 i_38_138 (.A1(n_449), .A2(n_75), .ZN(n_38_110));
   NAND2_X1 i_38_139 (.A1(n_450), .A2(n_74), .ZN(n_38_111));
   NAND2_X1 i_38_140 (.A1(n_452), .A2(multiplicand[27]), .ZN(n_38_112));
   NAND4_X1 i_38_141 (.A1(n_38_109), .A2(n_38_110), .A3(n_38_111), .A4(n_38_112), 
      .ZN(n_481));
   NAND2_X1 i_38_142 (.A1(n_451), .A2(multiplicand[29]), .ZN(n_38_113));
   NAND2_X1 i_38_143 (.A1(n_449), .A2(n_76), .ZN(n_38_114));
   NAND2_X1 i_38_144 (.A1(n_450), .A2(n_75), .ZN(n_38_115));
   NAND2_X1 i_38_145 (.A1(n_452), .A2(multiplicand[28]), .ZN(n_38_116));
   NAND4_X1 i_38_146 (.A1(n_38_113), .A2(n_38_114), .A3(n_38_115), .A4(n_38_116), 
      .ZN(n_482));
   NAND2_X1 i_38_147 (.A1(n_451), .A2(multiplicand[30]), .ZN(n_38_117));
   NAND2_X1 i_38_148 (.A1(n_449), .A2(n_77), .ZN(n_38_118));
   NAND2_X1 i_38_149 (.A1(n_450), .A2(n_76), .ZN(n_38_119));
   NAND2_X1 i_38_150 (.A1(n_452), .A2(multiplicand[29]), .ZN(n_38_120));
   NAND4_X1 i_38_151 (.A1(n_38_117), .A2(n_38_118), .A3(n_38_119), .A4(n_38_120), 
      .ZN(n_483));
   NAND2_X1 i_38_152 (.A1(n_451), .A2(multiplicand[31]), .ZN(n_38_121));
   NAND2_X1 i_38_153 (.A1(n_449), .A2(n_78), .ZN(n_38_122));
   NAND2_X1 i_38_154 (.A1(n_450), .A2(n_77), .ZN(n_38_123));
   NAND2_X1 i_38_155 (.A1(n_452), .A2(multiplicand[30]), .ZN(n_38_124));
   NAND4_X1 i_38_156 (.A1(n_38_121), .A2(n_38_122), .A3(n_38_123), .A4(n_38_124), 
      .ZN(n_484));
   NAND2_X1 i_38_157 (.A1(n_450), .A2(n_78), .ZN(n_38_125));
   NAND2_X1 i_38_158 (.A1(n_452), .A2(multiplicand[31]), .ZN(n_38_126));
   NAND4_X1 i_38_159 (.A1(n_38_121), .A2(n_38_122), .A3(n_38_125), .A4(n_38_126), 
      .ZN(n_485));
   INV_X1 i_39_0 (.A(n_33), .ZN(n_39_0));
   AND3_X1 i_39_1 (.A1(n_39_0), .A2(n_34), .A3(n_35), .ZN(n_486));
   INV_X1 i_39_2 (.A(n_34), .ZN(n_39_1));
   AND3_X1 i_39_3 (.A1(n_39_1), .A2(n_33), .A3(n_35), .ZN(n_487));
   NOR3_X1 i_39_4 (.A1(n_39_1), .A2(n_33), .A3(n_35), .ZN(n_488));
   NOR3_X1 i_39_5 (.A1(n_39_0), .A2(n_34), .A3(n_35), .ZN(n_489));
   AOI22_X1 i_40_0 (.A1(n_488), .A2(multiplicand[0]), .B1(n_486), .B2(
      multiplicand[0]), .ZN(n_40_0));
   INV_X1 i_40_1 (.A(n_40_0), .ZN(n_490));
   NAND2_X1 i_40_2 (.A1(n_488), .A2(multiplicand[1]), .ZN(n_40_1));
   NAND2_X1 i_40_3 (.A1(n_486), .A2(n_48), .ZN(n_40_2));
   NAND2_X1 i_40_4 (.A1(n_487), .A2(multiplicand[0]), .ZN(n_40_3));
   NAND2_X1 i_40_5 (.A1(n_489), .A2(multiplicand[0]), .ZN(n_40_4));
   NAND4_X1 i_40_6 (.A1(n_40_1), .A2(n_40_2), .A3(n_40_3), .A4(n_40_4), .ZN(
      n_491));
   NAND2_X1 i_40_7 (.A1(n_488), .A2(multiplicand[2]), .ZN(n_40_5));
   NAND2_X1 i_40_8 (.A1(n_486), .A2(n_49), .ZN(n_40_6));
   NAND2_X1 i_40_9 (.A1(n_487), .A2(n_48), .ZN(n_40_7));
   NAND2_X1 i_40_10 (.A1(n_489), .A2(multiplicand[1]), .ZN(n_40_8));
   NAND4_X1 i_40_11 (.A1(n_40_5), .A2(n_40_6), .A3(n_40_7), .A4(n_40_8), 
      .ZN(n_492));
   NAND2_X1 i_40_12 (.A1(n_488), .A2(multiplicand[3]), .ZN(n_40_9));
   NAND2_X1 i_40_13 (.A1(n_486), .A2(n_50), .ZN(n_40_10));
   NAND2_X1 i_40_14 (.A1(n_487), .A2(n_49), .ZN(n_40_11));
   NAND2_X1 i_40_15 (.A1(n_489), .A2(multiplicand[2]), .ZN(n_40_12));
   NAND4_X1 i_40_16 (.A1(n_40_9), .A2(n_40_10), .A3(n_40_11), .A4(n_40_12), 
      .ZN(n_493));
   NAND2_X1 i_40_17 (.A1(n_488), .A2(multiplicand[4]), .ZN(n_40_13));
   NAND2_X1 i_40_18 (.A1(n_486), .A2(n_51), .ZN(n_40_14));
   NAND2_X1 i_40_19 (.A1(n_487), .A2(n_50), .ZN(n_40_15));
   NAND2_X1 i_40_20 (.A1(n_489), .A2(multiplicand[3]), .ZN(n_40_16));
   NAND4_X1 i_40_21 (.A1(n_40_13), .A2(n_40_14), .A3(n_40_15), .A4(n_40_16), 
      .ZN(n_494));
   NAND2_X1 i_40_22 (.A1(n_488), .A2(multiplicand[5]), .ZN(n_40_17));
   NAND2_X1 i_40_23 (.A1(n_486), .A2(n_52), .ZN(n_40_18));
   NAND2_X1 i_40_24 (.A1(n_487), .A2(n_51), .ZN(n_40_19));
   NAND2_X1 i_40_25 (.A1(n_489), .A2(multiplicand[4]), .ZN(n_40_20));
   NAND4_X1 i_40_26 (.A1(n_40_17), .A2(n_40_18), .A3(n_40_19), .A4(n_40_20), 
      .ZN(n_495));
   NAND2_X1 i_40_27 (.A1(n_488), .A2(multiplicand[6]), .ZN(n_40_21));
   NAND2_X1 i_40_28 (.A1(n_486), .A2(n_53), .ZN(n_40_22));
   NAND2_X1 i_40_29 (.A1(n_487), .A2(n_52), .ZN(n_40_23));
   NAND2_X1 i_40_30 (.A1(n_489), .A2(multiplicand[5]), .ZN(n_40_24));
   NAND4_X1 i_40_31 (.A1(n_40_21), .A2(n_40_22), .A3(n_40_23), .A4(n_40_24), 
      .ZN(n_496));
   NAND2_X1 i_40_32 (.A1(n_488), .A2(multiplicand[7]), .ZN(n_40_25));
   NAND2_X1 i_40_33 (.A1(n_486), .A2(n_54), .ZN(n_40_26));
   NAND2_X1 i_40_34 (.A1(n_487), .A2(n_53), .ZN(n_40_27));
   NAND2_X1 i_40_35 (.A1(n_489), .A2(multiplicand[6]), .ZN(n_40_28));
   NAND4_X1 i_40_36 (.A1(n_40_25), .A2(n_40_26), .A3(n_40_27), .A4(n_40_28), 
      .ZN(n_497));
   NAND2_X1 i_40_37 (.A1(n_488), .A2(multiplicand[8]), .ZN(n_40_29));
   NAND2_X1 i_40_38 (.A1(n_486), .A2(n_55), .ZN(n_40_30));
   NAND2_X1 i_40_39 (.A1(n_487), .A2(n_54), .ZN(n_40_31));
   NAND2_X1 i_40_40 (.A1(n_489), .A2(multiplicand[7]), .ZN(n_40_32));
   NAND4_X1 i_40_41 (.A1(n_40_29), .A2(n_40_30), .A3(n_40_31), .A4(n_40_32), 
      .ZN(n_498));
   NAND2_X1 i_40_42 (.A1(n_488), .A2(multiplicand[9]), .ZN(n_40_33));
   NAND2_X1 i_40_43 (.A1(n_486), .A2(n_56), .ZN(n_40_34));
   NAND2_X1 i_40_44 (.A1(n_487), .A2(n_55), .ZN(n_40_35));
   NAND2_X1 i_40_45 (.A1(n_489), .A2(multiplicand[8]), .ZN(n_40_36));
   NAND4_X1 i_40_46 (.A1(n_40_33), .A2(n_40_34), .A3(n_40_35), .A4(n_40_36), 
      .ZN(n_499));
   NAND2_X1 i_40_47 (.A1(n_488), .A2(multiplicand[10]), .ZN(n_40_37));
   NAND2_X1 i_40_48 (.A1(n_486), .A2(n_57), .ZN(n_40_38));
   NAND2_X1 i_40_49 (.A1(n_487), .A2(n_56), .ZN(n_40_39));
   NAND2_X1 i_40_50 (.A1(n_489), .A2(multiplicand[9]), .ZN(n_40_40));
   NAND4_X1 i_40_51 (.A1(n_40_37), .A2(n_40_38), .A3(n_40_39), .A4(n_40_40), 
      .ZN(n_500));
   NAND2_X1 i_40_52 (.A1(n_488), .A2(multiplicand[11]), .ZN(n_40_41));
   NAND2_X1 i_40_53 (.A1(n_486), .A2(n_58), .ZN(n_40_42));
   NAND2_X1 i_40_54 (.A1(n_487), .A2(n_57), .ZN(n_40_43));
   NAND2_X1 i_40_55 (.A1(n_489), .A2(multiplicand[10]), .ZN(n_40_44));
   NAND4_X1 i_40_56 (.A1(n_40_41), .A2(n_40_42), .A3(n_40_43), .A4(n_40_44), 
      .ZN(n_501));
   NAND2_X1 i_40_57 (.A1(n_488), .A2(multiplicand[12]), .ZN(n_40_45));
   NAND2_X1 i_40_58 (.A1(n_486), .A2(n_59), .ZN(n_40_46));
   NAND2_X1 i_40_59 (.A1(n_487), .A2(n_58), .ZN(n_40_47));
   NAND2_X1 i_40_60 (.A1(n_489), .A2(multiplicand[11]), .ZN(n_40_48));
   NAND4_X1 i_40_61 (.A1(n_40_45), .A2(n_40_46), .A3(n_40_47), .A4(n_40_48), 
      .ZN(n_502));
   NAND2_X1 i_40_62 (.A1(n_488), .A2(multiplicand[13]), .ZN(n_40_49));
   NAND2_X1 i_40_63 (.A1(n_486), .A2(n_60), .ZN(n_40_50));
   NAND2_X1 i_40_64 (.A1(n_487), .A2(n_59), .ZN(n_40_51));
   NAND2_X1 i_40_65 (.A1(n_489), .A2(multiplicand[12]), .ZN(n_40_52));
   NAND4_X1 i_40_66 (.A1(n_40_49), .A2(n_40_50), .A3(n_40_51), .A4(n_40_52), 
      .ZN(n_503));
   NAND2_X1 i_40_67 (.A1(n_488), .A2(multiplicand[14]), .ZN(n_40_53));
   NAND2_X1 i_40_68 (.A1(n_486), .A2(n_61), .ZN(n_40_54));
   NAND2_X1 i_40_69 (.A1(n_487), .A2(n_60), .ZN(n_40_55));
   NAND2_X1 i_40_70 (.A1(n_489), .A2(multiplicand[13]), .ZN(n_40_56));
   NAND4_X1 i_40_71 (.A1(n_40_53), .A2(n_40_54), .A3(n_40_55), .A4(n_40_56), 
      .ZN(n_504));
   NAND2_X1 i_40_72 (.A1(n_488), .A2(multiplicand[15]), .ZN(n_40_57));
   NAND2_X1 i_40_73 (.A1(n_486), .A2(n_62), .ZN(n_40_58));
   NAND2_X1 i_40_74 (.A1(n_487), .A2(n_61), .ZN(n_40_59));
   NAND2_X1 i_40_75 (.A1(n_489), .A2(multiplicand[14]), .ZN(n_40_60));
   NAND4_X1 i_40_76 (.A1(n_40_57), .A2(n_40_58), .A3(n_40_59), .A4(n_40_60), 
      .ZN(n_505));
   NAND2_X1 i_40_77 (.A1(n_488), .A2(multiplicand[16]), .ZN(n_40_61));
   NAND2_X1 i_40_78 (.A1(n_486), .A2(n_63), .ZN(n_40_62));
   NAND2_X1 i_40_79 (.A1(n_487), .A2(n_62), .ZN(n_40_63));
   NAND2_X1 i_40_80 (.A1(n_489), .A2(multiplicand[15]), .ZN(n_40_64));
   NAND4_X1 i_40_81 (.A1(n_40_61), .A2(n_40_62), .A3(n_40_63), .A4(n_40_64), 
      .ZN(n_506));
   NAND2_X1 i_40_82 (.A1(n_488), .A2(multiplicand[17]), .ZN(n_40_65));
   NAND2_X1 i_40_83 (.A1(n_486), .A2(n_64), .ZN(n_40_66));
   NAND2_X1 i_40_84 (.A1(n_487), .A2(n_63), .ZN(n_40_67));
   NAND2_X1 i_40_85 (.A1(n_489), .A2(multiplicand[16]), .ZN(n_40_68));
   NAND4_X1 i_40_86 (.A1(n_40_65), .A2(n_40_66), .A3(n_40_67), .A4(n_40_68), 
      .ZN(n_507));
   NAND2_X1 i_40_87 (.A1(n_488), .A2(multiplicand[18]), .ZN(n_40_69));
   NAND2_X1 i_40_88 (.A1(n_486), .A2(n_65), .ZN(n_40_70));
   NAND2_X1 i_40_89 (.A1(n_487), .A2(n_64), .ZN(n_40_71));
   NAND2_X1 i_40_90 (.A1(n_489), .A2(multiplicand[17]), .ZN(n_40_72));
   NAND4_X1 i_40_91 (.A1(n_40_69), .A2(n_40_70), .A3(n_40_71), .A4(n_40_72), 
      .ZN(n_508));
   NAND2_X1 i_40_92 (.A1(n_488), .A2(multiplicand[19]), .ZN(n_40_73));
   NAND2_X1 i_40_93 (.A1(n_486), .A2(n_66), .ZN(n_40_74));
   NAND2_X1 i_40_94 (.A1(n_487), .A2(n_65), .ZN(n_40_75));
   NAND2_X1 i_40_95 (.A1(n_489), .A2(multiplicand[18]), .ZN(n_40_76));
   NAND4_X1 i_40_96 (.A1(n_40_73), .A2(n_40_74), .A3(n_40_75), .A4(n_40_76), 
      .ZN(n_509));
   NAND2_X1 i_40_97 (.A1(n_488), .A2(multiplicand[20]), .ZN(n_40_77));
   NAND2_X1 i_40_98 (.A1(n_486), .A2(n_67), .ZN(n_40_78));
   NAND2_X1 i_40_99 (.A1(n_487), .A2(n_66), .ZN(n_40_79));
   NAND2_X1 i_40_100 (.A1(n_489), .A2(multiplicand[19]), .ZN(n_40_80));
   NAND4_X1 i_40_101 (.A1(n_40_77), .A2(n_40_78), .A3(n_40_79), .A4(n_40_80), 
      .ZN(n_510));
   NAND2_X1 i_40_102 (.A1(n_488), .A2(multiplicand[21]), .ZN(n_40_81));
   NAND2_X1 i_40_103 (.A1(n_486), .A2(n_68), .ZN(n_40_82));
   NAND2_X1 i_40_104 (.A1(n_487), .A2(n_67), .ZN(n_40_83));
   NAND2_X1 i_40_105 (.A1(n_489), .A2(multiplicand[20]), .ZN(n_40_84));
   NAND4_X1 i_40_106 (.A1(n_40_81), .A2(n_40_82), .A3(n_40_83), .A4(n_40_84), 
      .ZN(n_511));
   NAND2_X1 i_40_107 (.A1(n_488), .A2(multiplicand[22]), .ZN(n_40_85));
   NAND2_X1 i_40_108 (.A1(n_486), .A2(n_69), .ZN(n_40_86));
   NAND2_X1 i_40_109 (.A1(n_487), .A2(n_68), .ZN(n_40_87));
   NAND2_X1 i_40_110 (.A1(n_489), .A2(multiplicand[21]), .ZN(n_40_88));
   NAND4_X1 i_40_111 (.A1(n_40_85), .A2(n_40_86), .A3(n_40_87), .A4(n_40_88), 
      .ZN(n_512));
   NAND2_X1 i_40_112 (.A1(n_488), .A2(multiplicand[23]), .ZN(n_40_89));
   NAND2_X1 i_40_113 (.A1(n_486), .A2(n_70), .ZN(n_40_90));
   NAND2_X1 i_40_114 (.A1(n_487), .A2(n_69), .ZN(n_40_91));
   NAND2_X1 i_40_115 (.A1(n_489), .A2(multiplicand[22]), .ZN(n_40_92));
   NAND4_X1 i_40_116 (.A1(n_40_89), .A2(n_40_90), .A3(n_40_91), .A4(n_40_92), 
      .ZN(n_513));
   NAND2_X1 i_40_117 (.A1(n_488), .A2(multiplicand[24]), .ZN(n_40_93));
   NAND2_X1 i_40_118 (.A1(n_486), .A2(n_71), .ZN(n_40_94));
   NAND2_X1 i_40_119 (.A1(n_487), .A2(n_70), .ZN(n_40_95));
   NAND2_X1 i_40_120 (.A1(n_489), .A2(multiplicand[23]), .ZN(n_40_96));
   NAND4_X1 i_40_121 (.A1(n_40_93), .A2(n_40_94), .A3(n_40_95), .A4(n_40_96), 
      .ZN(n_514));
   NAND2_X1 i_40_122 (.A1(n_488), .A2(multiplicand[25]), .ZN(n_40_97));
   NAND2_X1 i_40_123 (.A1(n_486), .A2(n_72), .ZN(n_40_98));
   NAND2_X1 i_40_124 (.A1(n_487), .A2(n_71), .ZN(n_40_99));
   NAND2_X1 i_40_125 (.A1(n_489), .A2(multiplicand[24]), .ZN(n_40_100));
   NAND4_X1 i_40_126 (.A1(n_40_97), .A2(n_40_98), .A3(n_40_99), .A4(n_40_100), 
      .ZN(n_515));
   NAND2_X1 i_40_127 (.A1(n_488), .A2(multiplicand[26]), .ZN(n_40_101));
   NAND2_X1 i_40_128 (.A1(n_486), .A2(n_73), .ZN(n_40_102));
   NAND2_X1 i_40_129 (.A1(n_487), .A2(n_72), .ZN(n_40_103));
   NAND2_X1 i_40_130 (.A1(n_489), .A2(multiplicand[25]), .ZN(n_40_104));
   NAND4_X1 i_40_131 (.A1(n_40_101), .A2(n_40_102), .A3(n_40_103), .A4(n_40_104), 
      .ZN(n_516));
   NAND2_X1 i_40_132 (.A1(n_488), .A2(multiplicand[27]), .ZN(n_40_105));
   NAND2_X1 i_40_133 (.A1(n_486), .A2(n_74), .ZN(n_40_106));
   NAND2_X1 i_40_134 (.A1(n_487), .A2(n_73), .ZN(n_40_107));
   NAND2_X1 i_40_135 (.A1(n_489), .A2(multiplicand[26]), .ZN(n_40_108));
   NAND4_X1 i_40_136 (.A1(n_40_105), .A2(n_40_106), .A3(n_40_107), .A4(n_40_108), 
      .ZN(n_517));
   NAND2_X1 i_40_137 (.A1(n_488), .A2(multiplicand[28]), .ZN(n_40_109));
   NAND2_X1 i_40_138 (.A1(n_486), .A2(n_75), .ZN(n_40_110));
   NAND2_X1 i_40_139 (.A1(n_487), .A2(n_74), .ZN(n_40_111));
   NAND2_X1 i_40_140 (.A1(n_489), .A2(multiplicand[27]), .ZN(n_40_112));
   NAND4_X1 i_40_141 (.A1(n_40_109), .A2(n_40_110), .A3(n_40_111), .A4(n_40_112), 
      .ZN(n_518));
   NAND2_X1 i_40_142 (.A1(n_488), .A2(multiplicand[29]), .ZN(n_40_113));
   NAND2_X1 i_40_143 (.A1(n_486), .A2(n_76), .ZN(n_40_114));
   NAND2_X1 i_40_144 (.A1(n_487), .A2(n_75), .ZN(n_40_115));
   NAND2_X1 i_40_145 (.A1(n_489), .A2(multiplicand[28]), .ZN(n_40_116));
   NAND4_X1 i_40_146 (.A1(n_40_113), .A2(n_40_114), .A3(n_40_115), .A4(n_40_116), 
      .ZN(n_519));
   NAND2_X1 i_40_147 (.A1(n_488), .A2(multiplicand[30]), .ZN(n_40_117));
   NAND2_X1 i_40_148 (.A1(n_486), .A2(n_77), .ZN(n_40_118));
   NAND2_X1 i_40_149 (.A1(n_487), .A2(n_76), .ZN(n_40_119));
   NAND2_X1 i_40_150 (.A1(n_489), .A2(multiplicand[29]), .ZN(n_40_120));
   NAND4_X1 i_40_151 (.A1(n_40_117), .A2(n_40_118), .A3(n_40_119), .A4(n_40_120), 
      .ZN(n_520));
   NAND2_X1 i_40_152 (.A1(n_488), .A2(multiplicand[31]), .ZN(n_40_121));
   NAND2_X1 i_40_153 (.A1(n_486), .A2(n_78), .ZN(n_40_122));
   NAND2_X1 i_40_154 (.A1(n_487), .A2(n_77), .ZN(n_40_123));
   NAND2_X1 i_40_155 (.A1(n_489), .A2(multiplicand[30]), .ZN(n_40_124));
   NAND4_X1 i_40_156 (.A1(n_40_121), .A2(n_40_122), .A3(n_40_123), .A4(n_40_124), 
      .ZN(n_521));
   NAND2_X1 i_40_157 (.A1(n_487), .A2(n_78), .ZN(n_40_125));
   NAND2_X1 i_40_158 (.A1(n_489), .A2(multiplicand[31]), .ZN(n_40_126));
   NAND4_X1 i_40_159 (.A1(n_40_121), .A2(n_40_122), .A3(n_40_125), .A4(n_40_126), 
      .ZN(n_522));
   INV_X1 i_41_0 (.A(n_36), .ZN(n_41_0));
   AND3_X1 i_41_1 (.A1(n_41_0), .A2(n_37), .A3(n_38), .ZN(n_523));
   INV_X1 i_41_2 (.A(n_37), .ZN(n_41_1));
   AND3_X1 i_41_3 (.A1(n_41_1), .A2(n_36), .A3(n_38), .ZN(n_524));
   NOR3_X1 i_41_4 (.A1(n_41_1), .A2(n_36), .A3(n_38), .ZN(n_525));
   NOR3_X1 i_41_5 (.A1(n_41_0), .A2(n_37), .A3(n_38), .ZN(n_526));
   AOI22_X1 i_42_0 (.A1(n_525), .A2(multiplicand[0]), .B1(n_523), .B2(
      multiplicand[0]), .ZN(n_42_0));
   INV_X1 i_42_1 (.A(n_42_0), .ZN(n_527));
   NAND2_X1 i_42_2 (.A1(n_525), .A2(multiplicand[1]), .ZN(n_42_1));
   NAND2_X1 i_42_3 (.A1(n_523), .A2(n_48), .ZN(n_42_2));
   NAND2_X1 i_42_4 (.A1(n_524), .A2(multiplicand[0]), .ZN(n_42_3));
   NAND2_X1 i_42_5 (.A1(n_526), .A2(multiplicand[0]), .ZN(n_42_4));
   NAND4_X1 i_42_6 (.A1(n_42_1), .A2(n_42_2), .A3(n_42_3), .A4(n_42_4), .ZN(
      n_528));
   NAND2_X1 i_42_7 (.A1(n_525), .A2(multiplicand[2]), .ZN(n_42_5));
   NAND2_X1 i_42_8 (.A1(n_523), .A2(n_49), .ZN(n_42_6));
   NAND2_X1 i_42_9 (.A1(n_524), .A2(n_48), .ZN(n_42_7));
   NAND2_X1 i_42_10 (.A1(n_526), .A2(multiplicand[1]), .ZN(n_42_8));
   NAND4_X1 i_42_11 (.A1(n_42_5), .A2(n_42_6), .A3(n_42_7), .A4(n_42_8), 
      .ZN(n_529));
   NAND2_X1 i_42_12 (.A1(n_525), .A2(multiplicand[3]), .ZN(n_42_9));
   NAND2_X1 i_42_13 (.A1(n_523), .A2(n_50), .ZN(n_42_10));
   NAND2_X1 i_42_14 (.A1(n_524), .A2(n_49), .ZN(n_42_11));
   NAND2_X1 i_42_15 (.A1(n_526), .A2(multiplicand[2]), .ZN(n_42_12));
   NAND4_X1 i_42_16 (.A1(n_42_9), .A2(n_42_10), .A3(n_42_11), .A4(n_42_12), 
      .ZN(n_530));
   NAND2_X1 i_42_17 (.A1(n_525), .A2(multiplicand[4]), .ZN(n_42_13));
   NAND2_X1 i_42_18 (.A1(n_523), .A2(n_51), .ZN(n_42_14));
   NAND2_X1 i_42_19 (.A1(n_524), .A2(n_50), .ZN(n_42_15));
   NAND2_X1 i_42_20 (.A1(n_526), .A2(multiplicand[3]), .ZN(n_42_16));
   NAND4_X1 i_42_21 (.A1(n_42_13), .A2(n_42_14), .A3(n_42_15), .A4(n_42_16), 
      .ZN(n_531));
   NAND2_X1 i_42_22 (.A1(n_525), .A2(multiplicand[5]), .ZN(n_42_17));
   NAND2_X1 i_42_23 (.A1(n_523), .A2(n_52), .ZN(n_42_18));
   NAND2_X1 i_42_24 (.A1(n_524), .A2(n_51), .ZN(n_42_19));
   NAND2_X1 i_42_25 (.A1(n_526), .A2(multiplicand[4]), .ZN(n_42_20));
   NAND4_X1 i_42_26 (.A1(n_42_17), .A2(n_42_18), .A3(n_42_19), .A4(n_42_20), 
      .ZN(n_532));
   NAND2_X1 i_42_27 (.A1(n_525), .A2(multiplicand[6]), .ZN(n_42_21));
   NAND2_X1 i_42_28 (.A1(n_523), .A2(n_53), .ZN(n_42_22));
   NAND2_X1 i_42_29 (.A1(n_524), .A2(n_52), .ZN(n_42_23));
   NAND2_X1 i_42_30 (.A1(n_526), .A2(multiplicand[5]), .ZN(n_42_24));
   NAND4_X1 i_42_31 (.A1(n_42_21), .A2(n_42_22), .A3(n_42_23), .A4(n_42_24), 
      .ZN(n_533));
   NAND2_X1 i_42_32 (.A1(n_525), .A2(multiplicand[7]), .ZN(n_42_25));
   NAND2_X1 i_42_33 (.A1(n_523), .A2(n_54), .ZN(n_42_26));
   NAND2_X1 i_42_34 (.A1(n_524), .A2(n_53), .ZN(n_42_27));
   NAND2_X1 i_42_35 (.A1(n_526), .A2(multiplicand[6]), .ZN(n_42_28));
   NAND4_X1 i_42_36 (.A1(n_42_25), .A2(n_42_26), .A3(n_42_27), .A4(n_42_28), 
      .ZN(n_534));
   NAND2_X1 i_42_37 (.A1(n_525), .A2(multiplicand[8]), .ZN(n_42_29));
   NAND2_X1 i_42_38 (.A1(n_523), .A2(n_55), .ZN(n_42_30));
   NAND2_X1 i_42_39 (.A1(n_524), .A2(n_54), .ZN(n_42_31));
   NAND2_X1 i_42_40 (.A1(n_526), .A2(multiplicand[7]), .ZN(n_42_32));
   NAND4_X1 i_42_41 (.A1(n_42_29), .A2(n_42_30), .A3(n_42_31), .A4(n_42_32), 
      .ZN(n_535));
   NAND2_X1 i_42_42 (.A1(n_525), .A2(multiplicand[9]), .ZN(n_42_33));
   NAND2_X1 i_42_43 (.A1(n_523), .A2(n_56), .ZN(n_42_34));
   NAND2_X1 i_42_44 (.A1(n_524), .A2(n_55), .ZN(n_42_35));
   NAND2_X1 i_42_45 (.A1(n_526), .A2(multiplicand[8]), .ZN(n_42_36));
   NAND4_X1 i_42_46 (.A1(n_42_33), .A2(n_42_34), .A3(n_42_35), .A4(n_42_36), 
      .ZN(n_536));
   NAND2_X1 i_42_47 (.A1(n_525), .A2(multiplicand[10]), .ZN(n_42_37));
   NAND2_X1 i_42_48 (.A1(n_523), .A2(n_57), .ZN(n_42_38));
   NAND2_X1 i_42_49 (.A1(n_524), .A2(n_56), .ZN(n_42_39));
   NAND2_X1 i_42_50 (.A1(n_526), .A2(multiplicand[9]), .ZN(n_42_40));
   NAND4_X1 i_42_51 (.A1(n_42_37), .A2(n_42_38), .A3(n_42_39), .A4(n_42_40), 
      .ZN(n_537));
   NAND2_X1 i_42_52 (.A1(n_525), .A2(multiplicand[11]), .ZN(n_42_41));
   NAND2_X1 i_42_53 (.A1(n_523), .A2(n_58), .ZN(n_42_42));
   NAND2_X1 i_42_54 (.A1(n_524), .A2(n_57), .ZN(n_42_43));
   NAND2_X1 i_42_55 (.A1(n_526), .A2(multiplicand[10]), .ZN(n_42_44));
   NAND4_X1 i_42_56 (.A1(n_42_41), .A2(n_42_42), .A3(n_42_43), .A4(n_42_44), 
      .ZN(n_538));
   NAND2_X1 i_42_57 (.A1(n_525), .A2(multiplicand[12]), .ZN(n_42_45));
   NAND2_X1 i_42_58 (.A1(n_523), .A2(n_59), .ZN(n_42_46));
   NAND2_X1 i_42_59 (.A1(n_524), .A2(n_58), .ZN(n_42_47));
   NAND2_X1 i_42_60 (.A1(n_526), .A2(multiplicand[11]), .ZN(n_42_48));
   NAND4_X1 i_42_61 (.A1(n_42_45), .A2(n_42_46), .A3(n_42_47), .A4(n_42_48), 
      .ZN(n_539));
   NAND2_X1 i_42_62 (.A1(n_525), .A2(multiplicand[13]), .ZN(n_42_49));
   NAND2_X1 i_42_63 (.A1(n_523), .A2(n_60), .ZN(n_42_50));
   NAND2_X1 i_42_64 (.A1(n_524), .A2(n_59), .ZN(n_42_51));
   NAND2_X1 i_42_65 (.A1(n_526), .A2(multiplicand[12]), .ZN(n_42_52));
   NAND4_X1 i_42_66 (.A1(n_42_49), .A2(n_42_50), .A3(n_42_51), .A4(n_42_52), 
      .ZN(n_540));
   NAND2_X1 i_42_67 (.A1(n_525), .A2(multiplicand[14]), .ZN(n_42_53));
   NAND2_X1 i_42_68 (.A1(n_523), .A2(n_61), .ZN(n_42_54));
   NAND2_X1 i_42_69 (.A1(n_524), .A2(n_60), .ZN(n_42_55));
   NAND2_X1 i_42_70 (.A1(n_526), .A2(multiplicand[13]), .ZN(n_42_56));
   NAND4_X1 i_42_71 (.A1(n_42_53), .A2(n_42_54), .A3(n_42_55), .A4(n_42_56), 
      .ZN(n_541));
   NAND2_X1 i_42_72 (.A1(n_525), .A2(multiplicand[15]), .ZN(n_42_57));
   NAND2_X1 i_42_73 (.A1(n_523), .A2(n_62), .ZN(n_42_58));
   NAND2_X1 i_42_74 (.A1(n_524), .A2(n_61), .ZN(n_42_59));
   NAND2_X1 i_42_75 (.A1(n_526), .A2(multiplicand[14]), .ZN(n_42_60));
   NAND4_X1 i_42_76 (.A1(n_42_57), .A2(n_42_58), .A3(n_42_59), .A4(n_42_60), 
      .ZN(n_542));
   NAND2_X1 i_42_77 (.A1(n_525), .A2(multiplicand[16]), .ZN(n_42_61));
   NAND2_X1 i_42_78 (.A1(n_523), .A2(n_63), .ZN(n_42_62));
   NAND2_X1 i_42_79 (.A1(n_524), .A2(n_62), .ZN(n_42_63));
   NAND2_X1 i_42_80 (.A1(n_526), .A2(multiplicand[15]), .ZN(n_42_64));
   NAND4_X1 i_42_81 (.A1(n_42_61), .A2(n_42_62), .A3(n_42_63), .A4(n_42_64), 
      .ZN(n_543));
   NAND2_X1 i_42_82 (.A1(n_525), .A2(multiplicand[17]), .ZN(n_42_65));
   NAND2_X1 i_42_83 (.A1(n_523), .A2(n_64), .ZN(n_42_66));
   NAND2_X1 i_42_84 (.A1(n_524), .A2(n_63), .ZN(n_42_67));
   NAND2_X1 i_42_85 (.A1(n_526), .A2(multiplicand[16]), .ZN(n_42_68));
   NAND4_X1 i_42_86 (.A1(n_42_65), .A2(n_42_66), .A3(n_42_67), .A4(n_42_68), 
      .ZN(n_544));
   NAND2_X1 i_42_87 (.A1(n_525), .A2(multiplicand[18]), .ZN(n_42_69));
   NAND2_X1 i_42_88 (.A1(n_523), .A2(n_65), .ZN(n_42_70));
   NAND2_X1 i_42_89 (.A1(n_524), .A2(n_64), .ZN(n_42_71));
   NAND2_X1 i_42_90 (.A1(n_526), .A2(multiplicand[17]), .ZN(n_42_72));
   NAND4_X1 i_42_91 (.A1(n_42_69), .A2(n_42_70), .A3(n_42_71), .A4(n_42_72), 
      .ZN(n_545));
   NAND2_X1 i_42_92 (.A1(n_525), .A2(multiplicand[19]), .ZN(n_42_73));
   NAND2_X1 i_42_93 (.A1(n_523), .A2(n_66), .ZN(n_42_74));
   NAND2_X1 i_42_94 (.A1(n_524), .A2(n_65), .ZN(n_42_75));
   NAND2_X1 i_42_95 (.A1(n_526), .A2(multiplicand[18]), .ZN(n_42_76));
   NAND4_X1 i_42_96 (.A1(n_42_73), .A2(n_42_74), .A3(n_42_75), .A4(n_42_76), 
      .ZN(n_546));
   NAND2_X1 i_42_97 (.A1(n_525), .A2(multiplicand[20]), .ZN(n_42_77));
   NAND2_X1 i_42_98 (.A1(n_523), .A2(n_67), .ZN(n_42_78));
   NAND2_X1 i_42_99 (.A1(n_524), .A2(n_66), .ZN(n_42_79));
   NAND2_X1 i_42_100 (.A1(n_526), .A2(multiplicand[19]), .ZN(n_42_80));
   NAND4_X1 i_42_101 (.A1(n_42_77), .A2(n_42_78), .A3(n_42_79), .A4(n_42_80), 
      .ZN(n_547));
   NAND2_X1 i_42_102 (.A1(n_525), .A2(multiplicand[21]), .ZN(n_42_81));
   NAND2_X1 i_42_103 (.A1(n_523), .A2(n_68), .ZN(n_42_82));
   NAND2_X1 i_42_104 (.A1(n_524), .A2(n_67), .ZN(n_42_83));
   NAND2_X1 i_42_105 (.A1(n_526), .A2(multiplicand[20]), .ZN(n_42_84));
   NAND4_X1 i_42_106 (.A1(n_42_81), .A2(n_42_82), .A3(n_42_83), .A4(n_42_84), 
      .ZN(n_548));
   NAND2_X1 i_42_107 (.A1(n_525), .A2(multiplicand[22]), .ZN(n_42_85));
   NAND2_X1 i_42_108 (.A1(n_523), .A2(n_69), .ZN(n_42_86));
   NAND2_X1 i_42_109 (.A1(n_524), .A2(n_68), .ZN(n_42_87));
   NAND2_X1 i_42_110 (.A1(n_526), .A2(multiplicand[21]), .ZN(n_42_88));
   NAND4_X1 i_42_111 (.A1(n_42_85), .A2(n_42_86), .A3(n_42_87), .A4(n_42_88), 
      .ZN(n_549));
   NAND2_X1 i_42_112 (.A1(n_525), .A2(multiplicand[23]), .ZN(n_42_89));
   NAND2_X1 i_42_113 (.A1(n_523), .A2(n_70), .ZN(n_42_90));
   NAND2_X1 i_42_114 (.A1(n_524), .A2(n_69), .ZN(n_42_91));
   NAND2_X1 i_42_115 (.A1(n_526), .A2(multiplicand[22]), .ZN(n_42_92));
   NAND4_X1 i_42_116 (.A1(n_42_89), .A2(n_42_90), .A3(n_42_91), .A4(n_42_92), 
      .ZN(n_550));
   NAND2_X1 i_42_117 (.A1(n_525), .A2(multiplicand[24]), .ZN(n_42_93));
   NAND2_X1 i_42_118 (.A1(n_523), .A2(n_71), .ZN(n_42_94));
   NAND2_X1 i_42_119 (.A1(n_524), .A2(n_70), .ZN(n_42_95));
   NAND2_X1 i_42_120 (.A1(n_526), .A2(multiplicand[23]), .ZN(n_42_96));
   NAND4_X1 i_42_121 (.A1(n_42_93), .A2(n_42_94), .A3(n_42_95), .A4(n_42_96), 
      .ZN(n_551));
   NAND2_X1 i_42_122 (.A1(n_525), .A2(multiplicand[25]), .ZN(n_42_97));
   NAND2_X1 i_42_123 (.A1(n_523), .A2(n_72), .ZN(n_42_98));
   NAND2_X1 i_42_124 (.A1(n_524), .A2(n_71), .ZN(n_42_99));
   NAND2_X1 i_42_125 (.A1(n_526), .A2(multiplicand[24]), .ZN(n_42_100));
   NAND4_X1 i_42_126 (.A1(n_42_97), .A2(n_42_98), .A3(n_42_99), .A4(n_42_100), 
      .ZN(n_552));
   NAND2_X1 i_42_127 (.A1(n_525), .A2(multiplicand[26]), .ZN(n_42_101));
   NAND2_X1 i_42_128 (.A1(n_523), .A2(n_73), .ZN(n_42_102));
   NAND2_X1 i_42_129 (.A1(n_524), .A2(n_72), .ZN(n_42_103));
   NAND2_X1 i_42_130 (.A1(n_526), .A2(multiplicand[25]), .ZN(n_42_104));
   NAND4_X1 i_42_131 (.A1(n_42_101), .A2(n_42_102), .A3(n_42_103), .A4(n_42_104), 
      .ZN(n_553));
   NAND2_X1 i_42_132 (.A1(n_525), .A2(multiplicand[27]), .ZN(n_42_105));
   NAND2_X1 i_42_133 (.A1(n_523), .A2(n_74), .ZN(n_42_106));
   NAND2_X1 i_42_134 (.A1(n_524), .A2(n_73), .ZN(n_42_107));
   NAND2_X1 i_42_135 (.A1(n_526), .A2(multiplicand[26]), .ZN(n_42_108));
   NAND4_X1 i_42_136 (.A1(n_42_105), .A2(n_42_106), .A3(n_42_107), .A4(n_42_108), 
      .ZN(n_554));
   NAND2_X1 i_42_137 (.A1(n_525), .A2(multiplicand[28]), .ZN(n_42_109));
   NAND2_X1 i_42_138 (.A1(n_523), .A2(n_75), .ZN(n_42_110));
   NAND2_X1 i_42_139 (.A1(n_524), .A2(n_74), .ZN(n_42_111));
   NAND2_X1 i_42_140 (.A1(n_526), .A2(multiplicand[27]), .ZN(n_42_112));
   NAND4_X1 i_42_141 (.A1(n_42_109), .A2(n_42_110), .A3(n_42_111), .A4(n_42_112), 
      .ZN(n_555));
   NAND2_X1 i_42_142 (.A1(n_525), .A2(multiplicand[29]), .ZN(n_42_113));
   NAND2_X1 i_42_143 (.A1(n_523), .A2(n_76), .ZN(n_42_114));
   NAND2_X1 i_42_144 (.A1(n_524), .A2(n_75), .ZN(n_42_115));
   NAND2_X1 i_42_145 (.A1(n_526), .A2(multiplicand[28]), .ZN(n_42_116));
   NAND4_X1 i_42_146 (.A1(n_42_113), .A2(n_42_114), .A3(n_42_115), .A4(n_42_116), 
      .ZN(n_556));
   NAND2_X1 i_42_147 (.A1(n_525), .A2(multiplicand[30]), .ZN(n_42_117));
   NAND2_X1 i_42_148 (.A1(n_523), .A2(n_77), .ZN(n_42_118));
   NAND2_X1 i_42_149 (.A1(n_524), .A2(n_76), .ZN(n_42_119));
   NAND2_X1 i_42_150 (.A1(n_526), .A2(multiplicand[29]), .ZN(n_42_120));
   NAND4_X1 i_42_151 (.A1(n_42_117), .A2(n_42_118), .A3(n_42_119), .A4(n_42_120), 
      .ZN(n_557));
   NAND2_X1 i_42_152 (.A1(n_525), .A2(multiplicand[31]), .ZN(n_42_121));
   NAND2_X1 i_42_153 (.A1(n_523), .A2(n_78), .ZN(n_42_122));
   NAND2_X1 i_42_154 (.A1(n_524), .A2(n_77), .ZN(n_42_123));
   NAND2_X1 i_42_155 (.A1(n_526), .A2(multiplicand[30]), .ZN(n_42_124));
   NAND4_X1 i_42_156 (.A1(n_42_121), .A2(n_42_122), .A3(n_42_123), .A4(n_42_124), 
      .ZN(n_558));
   NAND2_X1 i_42_157 (.A1(n_524), .A2(n_78), .ZN(n_42_125));
   NAND2_X1 i_42_158 (.A1(n_526), .A2(multiplicand[31]), .ZN(n_42_126));
   NAND4_X1 i_42_159 (.A1(n_42_121), .A2(n_42_122), .A3(n_42_125), .A4(n_42_126), 
      .ZN(n_559));
   INV_X1 i_43_0 (.A(n_39), .ZN(n_43_0));
   AND3_X1 i_43_1 (.A1(n_43_0), .A2(n_40), .A3(n_41), .ZN(n_560));
   INV_X1 i_43_2 (.A(n_40), .ZN(n_43_1));
   AND3_X1 i_43_3 (.A1(n_43_1), .A2(n_39), .A3(n_41), .ZN(n_561));
   NOR3_X1 i_43_4 (.A1(n_43_1), .A2(n_39), .A3(n_41), .ZN(n_562));
   NOR3_X1 i_43_5 (.A1(n_43_0), .A2(n_40), .A3(n_41), .ZN(n_563));
   AOI22_X1 i_44_0 (.A1(n_562), .A2(multiplicand[0]), .B1(n_560), .B2(
      multiplicand[0]), .ZN(n_44_0));
   INV_X1 i_44_1 (.A(n_44_0), .ZN(n_564));
   NAND2_X1 i_44_2 (.A1(n_562), .A2(multiplicand[1]), .ZN(n_44_1));
   NAND2_X1 i_44_3 (.A1(n_560), .A2(n_48), .ZN(n_44_2));
   NAND2_X1 i_44_4 (.A1(n_561), .A2(multiplicand[0]), .ZN(n_44_3));
   NAND2_X1 i_44_5 (.A1(n_563), .A2(multiplicand[0]), .ZN(n_44_4));
   NAND4_X1 i_44_6 (.A1(n_44_1), .A2(n_44_2), .A3(n_44_3), .A4(n_44_4), .ZN(
      n_565));
   NAND2_X1 i_44_7 (.A1(n_562), .A2(multiplicand[2]), .ZN(n_44_5));
   NAND2_X1 i_44_8 (.A1(n_560), .A2(n_49), .ZN(n_44_6));
   NAND2_X1 i_44_9 (.A1(n_561), .A2(n_48), .ZN(n_44_7));
   NAND2_X1 i_44_10 (.A1(n_563), .A2(multiplicand[1]), .ZN(n_44_8));
   NAND4_X1 i_44_11 (.A1(n_44_5), .A2(n_44_6), .A3(n_44_7), .A4(n_44_8), 
      .ZN(n_566));
   NAND2_X1 i_44_12 (.A1(n_562), .A2(multiplicand[3]), .ZN(n_44_9));
   NAND2_X1 i_44_13 (.A1(n_560), .A2(n_50), .ZN(n_44_10));
   NAND2_X1 i_44_14 (.A1(n_561), .A2(n_49), .ZN(n_44_11));
   NAND2_X1 i_44_15 (.A1(n_563), .A2(multiplicand[2]), .ZN(n_44_12));
   NAND4_X1 i_44_16 (.A1(n_44_9), .A2(n_44_10), .A3(n_44_11), .A4(n_44_12), 
      .ZN(n_567));
   NAND2_X1 i_44_17 (.A1(n_562), .A2(multiplicand[4]), .ZN(n_44_13));
   NAND2_X1 i_44_18 (.A1(n_560), .A2(n_51), .ZN(n_44_14));
   NAND2_X1 i_44_19 (.A1(n_561), .A2(n_50), .ZN(n_44_15));
   NAND2_X1 i_44_20 (.A1(n_563), .A2(multiplicand[3]), .ZN(n_44_16));
   NAND4_X1 i_44_21 (.A1(n_44_13), .A2(n_44_14), .A3(n_44_15), .A4(n_44_16), 
      .ZN(n_568));
   NAND2_X1 i_44_22 (.A1(n_562), .A2(multiplicand[5]), .ZN(n_44_17));
   NAND2_X1 i_44_23 (.A1(n_560), .A2(n_52), .ZN(n_44_18));
   NAND2_X1 i_44_24 (.A1(n_561), .A2(n_51), .ZN(n_44_19));
   NAND2_X1 i_44_25 (.A1(n_563), .A2(multiplicand[4]), .ZN(n_44_20));
   NAND4_X1 i_44_26 (.A1(n_44_17), .A2(n_44_18), .A3(n_44_19), .A4(n_44_20), 
      .ZN(n_569));
   NAND2_X1 i_44_27 (.A1(n_562), .A2(multiplicand[6]), .ZN(n_44_21));
   NAND2_X1 i_44_28 (.A1(n_560), .A2(n_53), .ZN(n_44_22));
   NAND2_X1 i_44_29 (.A1(n_561), .A2(n_52), .ZN(n_44_23));
   NAND2_X1 i_44_30 (.A1(n_563), .A2(multiplicand[5]), .ZN(n_44_24));
   NAND4_X1 i_44_31 (.A1(n_44_21), .A2(n_44_22), .A3(n_44_23), .A4(n_44_24), 
      .ZN(n_570));
   NAND2_X1 i_44_32 (.A1(n_562), .A2(multiplicand[7]), .ZN(n_44_25));
   NAND2_X1 i_44_33 (.A1(n_560), .A2(n_54), .ZN(n_44_26));
   NAND2_X1 i_44_34 (.A1(n_561), .A2(n_53), .ZN(n_44_27));
   NAND2_X1 i_44_35 (.A1(n_563), .A2(multiplicand[6]), .ZN(n_44_28));
   NAND4_X1 i_44_36 (.A1(n_44_25), .A2(n_44_26), .A3(n_44_27), .A4(n_44_28), 
      .ZN(n_571));
   NAND2_X1 i_44_37 (.A1(n_562), .A2(multiplicand[8]), .ZN(n_44_29));
   NAND2_X1 i_44_38 (.A1(n_560), .A2(n_55), .ZN(n_44_30));
   NAND2_X1 i_44_39 (.A1(n_561), .A2(n_54), .ZN(n_44_31));
   NAND2_X1 i_44_40 (.A1(n_563), .A2(multiplicand[7]), .ZN(n_44_32));
   NAND4_X1 i_44_41 (.A1(n_44_29), .A2(n_44_30), .A3(n_44_31), .A4(n_44_32), 
      .ZN(n_572));
   NAND2_X1 i_44_42 (.A1(n_562), .A2(multiplicand[9]), .ZN(n_44_33));
   NAND2_X1 i_44_43 (.A1(n_560), .A2(n_56), .ZN(n_44_34));
   NAND2_X1 i_44_44 (.A1(n_561), .A2(n_55), .ZN(n_44_35));
   NAND2_X1 i_44_45 (.A1(n_563), .A2(multiplicand[8]), .ZN(n_44_36));
   NAND4_X1 i_44_46 (.A1(n_44_33), .A2(n_44_34), .A3(n_44_35), .A4(n_44_36), 
      .ZN(n_573));
   NAND2_X1 i_44_47 (.A1(n_562), .A2(multiplicand[10]), .ZN(n_44_37));
   NAND2_X1 i_44_48 (.A1(n_560), .A2(n_57), .ZN(n_44_38));
   NAND2_X1 i_44_49 (.A1(n_561), .A2(n_56), .ZN(n_44_39));
   NAND2_X1 i_44_50 (.A1(n_563), .A2(multiplicand[9]), .ZN(n_44_40));
   NAND4_X1 i_44_51 (.A1(n_44_37), .A2(n_44_38), .A3(n_44_39), .A4(n_44_40), 
      .ZN(n_574));
   NAND2_X1 i_44_52 (.A1(n_562), .A2(multiplicand[11]), .ZN(n_44_41));
   NAND2_X1 i_44_53 (.A1(n_560), .A2(n_58), .ZN(n_44_42));
   NAND2_X1 i_44_54 (.A1(n_561), .A2(n_57), .ZN(n_44_43));
   NAND2_X1 i_44_55 (.A1(n_563), .A2(multiplicand[10]), .ZN(n_44_44));
   NAND4_X1 i_44_56 (.A1(n_44_41), .A2(n_44_42), .A3(n_44_43), .A4(n_44_44), 
      .ZN(n_575));
   NAND2_X1 i_44_57 (.A1(n_562), .A2(multiplicand[12]), .ZN(n_44_45));
   NAND2_X1 i_44_58 (.A1(n_560), .A2(n_59), .ZN(n_44_46));
   NAND2_X1 i_44_59 (.A1(n_561), .A2(n_58), .ZN(n_44_47));
   NAND2_X1 i_44_60 (.A1(n_563), .A2(multiplicand[11]), .ZN(n_44_48));
   NAND4_X1 i_44_61 (.A1(n_44_45), .A2(n_44_46), .A3(n_44_47), .A4(n_44_48), 
      .ZN(n_576));
   NAND2_X1 i_44_62 (.A1(n_562), .A2(multiplicand[13]), .ZN(n_44_49));
   NAND2_X1 i_44_63 (.A1(n_560), .A2(n_60), .ZN(n_44_50));
   NAND2_X1 i_44_64 (.A1(n_561), .A2(n_59), .ZN(n_44_51));
   NAND2_X1 i_44_65 (.A1(n_563), .A2(multiplicand[12]), .ZN(n_44_52));
   NAND4_X1 i_44_66 (.A1(n_44_49), .A2(n_44_50), .A3(n_44_51), .A4(n_44_52), 
      .ZN(n_577));
   NAND2_X1 i_44_67 (.A1(n_562), .A2(multiplicand[14]), .ZN(n_44_53));
   NAND2_X1 i_44_68 (.A1(n_560), .A2(n_61), .ZN(n_44_54));
   NAND2_X1 i_44_69 (.A1(n_561), .A2(n_60), .ZN(n_44_55));
   NAND2_X1 i_44_70 (.A1(n_563), .A2(multiplicand[13]), .ZN(n_44_56));
   NAND4_X1 i_44_71 (.A1(n_44_53), .A2(n_44_54), .A3(n_44_55), .A4(n_44_56), 
      .ZN(n_578));
   NAND2_X1 i_44_72 (.A1(n_562), .A2(multiplicand[15]), .ZN(n_44_57));
   NAND2_X1 i_44_73 (.A1(n_560), .A2(n_62), .ZN(n_44_58));
   NAND2_X1 i_44_74 (.A1(n_561), .A2(n_61), .ZN(n_44_59));
   NAND2_X1 i_44_75 (.A1(n_563), .A2(multiplicand[14]), .ZN(n_44_60));
   NAND4_X1 i_44_76 (.A1(n_44_57), .A2(n_44_58), .A3(n_44_59), .A4(n_44_60), 
      .ZN(n_579));
   NAND2_X1 i_44_77 (.A1(n_562), .A2(multiplicand[16]), .ZN(n_44_61));
   NAND2_X1 i_44_78 (.A1(n_560), .A2(n_63), .ZN(n_44_62));
   NAND2_X1 i_44_79 (.A1(n_561), .A2(n_62), .ZN(n_44_63));
   NAND2_X1 i_44_80 (.A1(n_563), .A2(multiplicand[15]), .ZN(n_44_64));
   NAND4_X1 i_44_81 (.A1(n_44_61), .A2(n_44_62), .A3(n_44_63), .A4(n_44_64), 
      .ZN(n_580));
   NAND2_X1 i_44_82 (.A1(n_562), .A2(multiplicand[17]), .ZN(n_44_65));
   NAND2_X1 i_44_83 (.A1(n_560), .A2(n_64), .ZN(n_44_66));
   NAND2_X1 i_44_84 (.A1(n_561), .A2(n_63), .ZN(n_44_67));
   NAND2_X1 i_44_85 (.A1(n_563), .A2(multiplicand[16]), .ZN(n_44_68));
   NAND4_X1 i_44_86 (.A1(n_44_65), .A2(n_44_66), .A3(n_44_67), .A4(n_44_68), 
      .ZN(n_581));
   NAND2_X1 i_44_87 (.A1(n_562), .A2(multiplicand[18]), .ZN(n_44_69));
   NAND2_X1 i_44_88 (.A1(n_560), .A2(n_65), .ZN(n_44_70));
   NAND2_X1 i_44_89 (.A1(n_561), .A2(n_64), .ZN(n_44_71));
   NAND2_X1 i_44_90 (.A1(n_563), .A2(multiplicand[17]), .ZN(n_44_72));
   NAND4_X1 i_44_91 (.A1(n_44_69), .A2(n_44_70), .A3(n_44_71), .A4(n_44_72), 
      .ZN(n_582));
   NAND2_X1 i_44_92 (.A1(n_562), .A2(multiplicand[19]), .ZN(n_44_73));
   NAND2_X1 i_44_93 (.A1(n_560), .A2(n_66), .ZN(n_44_74));
   NAND2_X1 i_44_94 (.A1(n_561), .A2(n_65), .ZN(n_44_75));
   NAND2_X1 i_44_95 (.A1(n_563), .A2(multiplicand[18]), .ZN(n_44_76));
   NAND4_X1 i_44_96 (.A1(n_44_73), .A2(n_44_74), .A3(n_44_75), .A4(n_44_76), 
      .ZN(n_583));
   NAND2_X1 i_44_97 (.A1(n_562), .A2(multiplicand[20]), .ZN(n_44_77));
   NAND2_X1 i_44_98 (.A1(n_560), .A2(n_67), .ZN(n_44_78));
   NAND2_X1 i_44_99 (.A1(n_561), .A2(n_66), .ZN(n_44_79));
   NAND2_X1 i_44_100 (.A1(n_563), .A2(multiplicand[19]), .ZN(n_44_80));
   NAND4_X1 i_44_101 (.A1(n_44_77), .A2(n_44_78), .A3(n_44_79), .A4(n_44_80), 
      .ZN(n_584));
   NAND2_X1 i_44_102 (.A1(n_562), .A2(multiplicand[21]), .ZN(n_44_81));
   NAND2_X1 i_44_103 (.A1(n_560), .A2(n_68), .ZN(n_44_82));
   NAND2_X1 i_44_104 (.A1(n_561), .A2(n_67), .ZN(n_44_83));
   NAND2_X1 i_44_105 (.A1(n_563), .A2(multiplicand[20]), .ZN(n_44_84));
   NAND4_X1 i_44_106 (.A1(n_44_81), .A2(n_44_82), .A3(n_44_83), .A4(n_44_84), 
      .ZN(n_585));
   NAND2_X1 i_44_107 (.A1(n_562), .A2(multiplicand[22]), .ZN(n_44_85));
   NAND2_X1 i_44_108 (.A1(n_560), .A2(n_69), .ZN(n_44_86));
   NAND2_X1 i_44_109 (.A1(n_561), .A2(n_68), .ZN(n_44_87));
   NAND2_X1 i_44_110 (.A1(n_563), .A2(multiplicand[21]), .ZN(n_44_88));
   NAND4_X1 i_44_111 (.A1(n_44_85), .A2(n_44_86), .A3(n_44_87), .A4(n_44_88), 
      .ZN(n_586));
   NAND2_X1 i_44_112 (.A1(n_562), .A2(multiplicand[23]), .ZN(n_44_89));
   NAND2_X1 i_44_113 (.A1(n_560), .A2(n_70), .ZN(n_44_90));
   NAND2_X1 i_44_114 (.A1(n_561), .A2(n_69), .ZN(n_44_91));
   NAND2_X1 i_44_115 (.A1(n_563), .A2(multiplicand[22]), .ZN(n_44_92));
   NAND4_X1 i_44_116 (.A1(n_44_89), .A2(n_44_90), .A3(n_44_91), .A4(n_44_92), 
      .ZN(n_587));
   NAND2_X1 i_44_117 (.A1(n_562), .A2(multiplicand[24]), .ZN(n_44_93));
   NAND2_X1 i_44_118 (.A1(n_560), .A2(n_71), .ZN(n_44_94));
   NAND2_X1 i_44_119 (.A1(n_561), .A2(n_70), .ZN(n_44_95));
   NAND2_X1 i_44_120 (.A1(n_563), .A2(multiplicand[23]), .ZN(n_44_96));
   NAND4_X1 i_44_121 (.A1(n_44_93), .A2(n_44_94), .A3(n_44_95), .A4(n_44_96), 
      .ZN(n_588));
   NAND2_X1 i_44_122 (.A1(n_562), .A2(multiplicand[25]), .ZN(n_44_97));
   NAND2_X1 i_44_123 (.A1(n_560), .A2(n_72), .ZN(n_44_98));
   NAND2_X1 i_44_124 (.A1(n_561), .A2(n_71), .ZN(n_44_99));
   NAND2_X1 i_44_125 (.A1(n_563), .A2(multiplicand[24]), .ZN(n_44_100));
   NAND4_X1 i_44_126 (.A1(n_44_97), .A2(n_44_98), .A3(n_44_99), .A4(n_44_100), 
      .ZN(n_589));
   NAND2_X1 i_44_127 (.A1(n_562), .A2(multiplicand[26]), .ZN(n_44_101));
   NAND2_X1 i_44_128 (.A1(n_560), .A2(n_73), .ZN(n_44_102));
   NAND2_X1 i_44_129 (.A1(n_561), .A2(n_72), .ZN(n_44_103));
   NAND2_X1 i_44_130 (.A1(n_563), .A2(multiplicand[25]), .ZN(n_44_104));
   NAND4_X1 i_44_131 (.A1(n_44_101), .A2(n_44_102), .A3(n_44_103), .A4(n_44_104), 
      .ZN(n_590));
   NAND2_X1 i_44_132 (.A1(n_562), .A2(multiplicand[27]), .ZN(n_44_105));
   NAND2_X1 i_44_133 (.A1(n_560), .A2(n_74), .ZN(n_44_106));
   NAND2_X1 i_44_134 (.A1(n_561), .A2(n_73), .ZN(n_44_107));
   NAND2_X1 i_44_135 (.A1(n_563), .A2(multiplicand[26]), .ZN(n_44_108));
   NAND4_X1 i_44_136 (.A1(n_44_105), .A2(n_44_106), .A3(n_44_107), .A4(n_44_108), 
      .ZN(n_591));
   NAND2_X1 i_44_137 (.A1(n_562), .A2(multiplicand[28]), .ZN(n_44_109));
   NAND2_X1 i_44_138 (.A1(n_560), .A2(n_75), .ZN(n_44_110));
   NAND2_X1 i_44_139 (.A1(n_561), .A2(n_74), .ZN(n_44_111));
   NAND2_X1 i_44_140 (.A1(n_563), .A2(multiplicand[27]), .ZN(n_44_112));
   NAND4_X1 i_44_141 (.A1(n_44_109), .A2(n_44_110), .A3(n_44_111), .A4(n_44_112), 
      .ZN(n_592));
   NAND2_X1 i_44_142 (.A1(n_562), .A2(multiplicand[29]), .ZN(n_44_113));
   NAND2_X1 i_44_143 (.A1(n_560), .A2(n_76), .ZN(n_44_114));
   NAND2_X1 i_44_144 (.A1(n_561), .A2(n_75), .ZN(n_44_115));
   NAND2_X1 i_44_145 (.A1(n_563), .A2(multiplicand[28]), .ZN(n_44_116));
   NAND4_X1 i_44_146 (.A1(n_44_113), .A2(n_44_114), .A3(n_44_115), .A4(n_44_116), 
      .ZN(n_593));
   NAND2_X1 i_44_147 (.A1(n_562), .A2(multiplicand[30]), .ZN(n_44_117));
   NAND2_X1 i_44_148 (.A1(n_560), .A2(n_77), .ZN(n_44_118));
   NAND2_X1 i_44_149 (.A1(n_561), .A2(n_76), .ZN(n_44_119));
   NAND2_X1 i_44_150 (.A1(n_563), .A2(multiplicand[29]), .ZN(n_44_120));
   NAND4_X1 i_44_151 (.A1(n_44_117), .A2(n_44_118), .A3(n_44_119), .A4(n_44_120), 
      .ZN(n_594));
   NAND2_X1 i_44_152 (.A1(n_562), .A2(multiplicand[31]), .ZN(n_44_121));
   NAND2_X1 i_44_153 (.A1(n_560), .A2(n_78), .ZN(n_44_122));
   NAND2_X1 i_44_154 (.A1(n_561), .A2(n_77), .ZN(n_44_123));
   NAND2_X1 i_44_155 (.A1(n_563), .A2(multiplicand[30]), .ZN(n_44_124));
   NAND4_X1 i_44_156 (.A1(n_44_121), .A2(n_44_122), .A3(n_44_123), .A4(n_44_124), 
      .ZN(n_595));
   NAND2_X1 i_44_157 (.A1(n_561), .A2(n_78), .ZN(n_44_125));
   NAND2_X1 i_44_158 (.A1(n_563), .A2(multiplicand[31]), .ZN(n_44_126));
   NAND4_X1 i_44_159 (.A1(n_44_121), .A2(n_44_122), .A3(n_44_125), .A4(n_44_126), 
      .ZN(n_596));
   INV_X1 i_45_0 (.A(n_42), .ZN(n_45_0));
   AND3_X1 i_45_1 (.A1(n_45_0), .A2(n_43), .A3(n_44), .ZN(n_597));
   INV_X1 i_45_2 (.A(n_43), .ZN(n_45_1));
   AND3_X1 i_45_3 (.A1(n_45_1), .A2(n_42), .A3(n_44), .ZN(n_598));
   NOR3_X1 i_45_4 (.A1(n_45_1), .A2(n_42), .A3(n_44), .ZN(n_599));
   NOR3_X1 i_45_5 (.A1(n_45_0), .A2(n_43), .A3(n_44), .ZN(n_600));
   AOI22_X1 i_46_0 (.A1(n_599), .A2(multiplicand[0]), .B1(n_597), .B2(
      multiplicand[0]), .ZN(n_46_0));
   INV_X1 i_46_1 (.A(n_46_0), .ZN(n_601));
   NAND2_X1 i_46_2 (.A1(n_599), .A2(multiplicand[1]), .ZN(n_46_1));
   NAND2_X1 i_46_3 (.A1(n_597), .A2(n_48), .ZN(n_46_2));
   NAND2_X1 i_46_4 (.A1(n_598), .A2(multiplicand[0]), .ZN(n_46_3));
   NAND2_X1 i_46_5 (.A1(n_600), .A2(multiplicand[0]), .ZN(n_46_4));
   NAND4_X1 i_46_6 (.A1(n_46_1), .A2(n_46_2), .A3(n_46_3), .A4(n_46_4), .ZN(
      n_602));
   NAND2_X1 i_46_7 (.A1(n_599), .A2(multiplicand[2]), .ZN(n_46_5));
   NAND2_X1 i_46_8 (.A1(n_597), .A2(n_49), .ZN(n_46_6));
   NAND2_X1 i_46_9 (.A1(n_598), .A2(n_48), .ZN(n_46_7));
   NAND2_X1 i_46_10 (.A1(n_600), .A2(multiplicand[1]), .ZN(n_46_8));
   NAND4_X1 i_46_11 (.A1(n_46_5), .A2(n_46_6), .A3(n_46_7), .A4(n_46_8), 
      .ZN(n_603));
   NAND2_X1 i_46_12 (.A1(n_599), .A2(multiplicand[3]), .ZN(n_46_9));
   NAND2_X1 i_46_13 (.A1(n_597), .A2(n_50), .ZN(n_46_10));
   NAND2_X1 i_46_14 (.A1(n_598), .A2(n_49), .ZN(n_46_11));
   NAND2_X1 i_46_15 (.A1(n_600), .A2(multiplicand[2]), .ZN(n_46_12));
   NAND4_X1 i_46_16 (.A1(n_46_9), .A2(n_46_10), .A3(n_46_11), .A4(n_46_12), 
      .ZN(n_604));
   NAND2_X1 i_46_17 (.A1(n_599), .A2(multiplicand[4]), .ZN(n_46_13));
   NAND2_X1 i_46_18 (.A1(n_597), .A2(n_51), .ZN(n_46_14));
   NAND2_X1 i_46_19 (.A1(n_598), .A2(n_50), .ZN(n_46_15));
   NAND2_X1 i_46_20 (.A1(n_600), .A2(multiplicand[3]), .ZN(n_46_16));
   NAND4_X1 i_46_21 (.A1(n_46_13), .A2(n_46_14), .A3(n_46_15), .A4(n_46_16), 
      .ZN(n_605));
   NAND2_X1 i_46_22 (.A1(n_599), .A2(multiplicand[5]), .ZN(n_46_17));
   NAND2_X1 i_46_23 (.A1(n_597), .A2(n_52), .ZN(n_46_18));
   NAND2_X1 i_46_24 (.A1(n_598), .A2(n_51), .ZN(n_46_19));
   NAND2_X1 i_46_25 (.A1(n_600), .A2(multiplicand[4]), .ZN(n_46_20));
   NAND4_X1 i_46_26 (.A1(n_46_17), .A2(n_46_18), .A3(n_46_19), .A4(n_46_20), 
      .ZN(n_606));
   NAND2_X1 i_46_27 (.A1(n_599), .A2(multiplicand[6]), .ZN(n_46_21));
   NAND2_X1 i_46_28 (.A1(n_597), .A2(n_53), .ZN(n_46_22));
   NAND2_X1 i_46_29 (.A1(n_598), .A2(n_52), .ZN(n_46_23));
   NAND2_X1 i_46_30 (.A1(n_600), .A2(multiplicand[5]), .ZN(n_46_24));
   NAND4_X1 i_46_31 (.A1(n_46_21), .A2(n_46_22), .A3(n_46_23), .A4(n_46_24), 
      .ZN(n_607));
   NAND2_X1 i_46_32 (.A1(n_599), .A2(multiplicand[7]), .ZN(n_46_25));
   NAND2_X1 i_46_33 (.A1(n_597), .A2(n_54), .ZN(n_46_26));
   NAND2_X1 i_46_34 (.A1(n_598), .A2(n_53), .ZN(n_46_27));
   NAND2_X1 i_46_35 (.A1(n_600), .A2(multiplicand[6]), .ZN(n_46_28));
   NAND4_X1 i_46_36 (.A1(n_46_25), .A2(n_46_26), .A3(n_46_27), .A4(n_46_28), 
      .ZN(n_608));
   NAND2_X1 i_46_37 (.A1(n_599), .A2(multiplicand[8]), .ZN(n_46_29));
   NAND2_X1 i_46_38 (.A1(n_597), .A2(n_55), .ZN(n_46_30));
   NAND2_X1 i_46_39 (.A1(n_598), .A2(n_54), .ZN(n_46_31));
   NAND2_X1 i_46_40 (.A1(n_600), .A2(multiplicand[7]), .ZN(n_46_32));
   NAND4_X1 i_46_41 (.A1(n_46_29), .A2(n_46_30), .A3(n_46_31), .A4(n_46_32), 
      .ZN(n_609));
   NAND2_X1 i_46_42 (.A1(n_599), .A2(multiplicand[9]), .ZN(n_46_33));
   NAND2_X1 i_46_43 (.A1(n_597), .A2(n_56), .ZN(n_46_34));
   NAND2_X1 i_46_44 (.A1(n_598), .A2(n_55), .ZN(n_46_35));
   NAND2_X1 i_46_45 (.A1(n_600), .A2(multiplicand[8]), .ZN(n_46_36));
   NAND4_X1 i_46_46 (.A1(n_46_33), .A2(n_46_34), .A3(n_46_35), .A4(n_46_36), 
      .ZN(n_610));
   NAND2_X1 i_46_47 (.A1(n_599), .A2(multiplicand[10]), .ZN(n_46_37));
   NAND2_X1 i_46_48 (.A1(n_597), .A2(n_57), .ZN(n_46_38));
   NAND2_X1 i_46_49 (.A1(n_598), .A2(n_56), .ZN(n_46_39));
   NAND2_X1 i_46_50 (.A1(n_600), .A2(multiplicand[9]), .ZN(n_46_40));
   NAND4_X1 i_46_51 (.A1(n_46_37), .A2(n_46_38), .A3(n_46_39), .A4(n_46_40), 
      .ZN(n_611));
   NAND2_X1 i_46_52 (.A1(n_599), .A2(multiplicand[11]), .ZN(n_46_41));
   NAND2_X1 i_46_53 (.A1(n_597), .A2(n_58), .ZN(n_46_42));
   NAND2_X1 i_46_54 (.A1(n_598), .A2(n_57), .ZN(n_46_43));
   NAND2_X1 i_46_55 (.A1(n_600), .A2(multiplicand[10]), .ZN(n_46_44));
   NAND4_X1 i_46_56 (.A1(n_46_41), .A2(n_46_42), .A3(n_46_43), .A4(n_46_44), 
      .ZN(n_612));
   NAND2_X1 i_46_57 (.A1(n_599), .A2(multiplicand[12]), .ZN(n_46_45));
   NAND2_X1 i_46_58 (.A1(n_597), .A2(n_59), .ZN(n_46_46));
   NAND2_X1 i_46_59 (.A1(n_598), .A2(n_58), .ZN(n_46_47));
   NAND2_X1 i_46_60 (.A1(n_600), .A2(multiplicand[11]), .ZN(n_46_48));
   NAND4_X1 i_46_61 (.A1(n_46_45), .A2(n_46_46), .A3(n_46_47), .A4(n_46_48), 
      .ZN(n_613));
   NAND2_X1 i_46_62 (.A1(n_599), .A2(multiplicand[13]), .ZN(n_46_49));
   NAND2_X1 i_46_63 (.A1(n_597), .A2(n_60), .ZN(n_46_50));
   NAND2_X1 i_46_64 (.A1(n_598), .A2(n_59), .ZN(n_46_51));
   NAND2_X1 i_46_65 (.A1(n_600), .A2(multiplicand[12]), .ZN(n_46_52));
   NAND4_X1 i_46_66 (.A1(n_46_49), .A2(n_46_50), .A3(n_46_51), .A4(n_46_52), 
      .ZN(n_614));
   NAND2_X1 i_46_67 (.A1(n_599), .A2(multiplicand[14]), .ZN(n_46_53));
   NAND2_X1 i_46_68 (.A1(n_597), .A2(n_61), .ZN(n_46_54));
   NAND2_X1 i_46_69 (.A1(n_598), .A2(n_60), .ZN(n_46_55));
   NAND2_X1 i_46_70 (.A1(n_600), .A2(multiplicand[13]), .ZN(n_46_56));
   NAND4_X1 i_46_71 (.A1(n_46_53), .A2(n_46_54), .A3(n_46_55), .A4(n_46_56), 
      .ZN(n_615));
   NAND2_X1 i_46_72 (.A1(n_599), .A2(multiplicand[15]), .ZN(n_46_57));
   NAND2_X1 i_46_73 (.A1(n_597), .A2(n_62), .ZN(n_46_58));
   NAND2_X1 i_46_74 (.A1(n_598), .A2(n_61), .ZN(n_46_59));
   NAND2_X1 i_46_75 (.A1(n_600), .A2(multiplicand[14]), .ZN(n_46_60));
   NAND4_X1 i_46_76 (.A1(n_46_57), .A2(n_46_58), .A3(n_46_59), .A4(n_46_60), 
      .ZN(n_616));
   NAND2_X1 i_46_77 (.A1(n_599), .A2(multiplicand[16]), .ZN(n_46_61));
   NAND2_X1 i_46_78 (.A1(n_597), .A2(n_63), .ZN(n_46_62));
   NAND2_X1 i_46_79 (.A1(n_598), .A2(n_62), .ZN(n_46_63));
   NAND2_X1 i_46_80 (.A1(n_600), .A2(multiplicand[15]), .ZN(n_46_64));
   NAND4_X1 i_46_81 (.A1(n_46_61), .A2(n_46_62), .A3(n_46_63), .A4(n_46_64), 
      .ZN(n_617));
   NAND2_X1 i_46_82 (.A1(n_599), .A2(multiplicand[17]), .ZN(n_46_65));
   NAND2_X1 i_46_83 (.A1(n_597), .A2(n_64), .ZN(n_46_66));
   NAND2_X1 i_46_84 (.A1(n_598), .A2(n_63), .ZN(n_46_67));
   NAND2_X1 i_46_85 (.A1(n_600), .A2(multiplicand[16]), .ZN(n_46_68));
   NAND4_X1 i_46_86 (.A1(n_46_65), .A2(n_46_66), .A3(n_46_67), .A4(n_46_68), 
      .ZN(n_618));
   NAND2_X1 i_46_87 (.A1(n_599), .A2(multiplicand[18]), .ZN(n_46_69));
   NAND2_X1 i_46_88 (.A1(n_597), .A2(n_65), .ZN(n_46_70));
   NAND2_X1 i_46_89 (.A1(n_598), .A2(n_64), .ZN(n_46_71));
   NAND2_X1 i_46_90 (.A1(n_600), .A2(multiplicand[17]), .ZN(n_46_72));
   NAND4_X1 i_46_91 (.A1(n_46_69), .A2(n_46_70), .A3(n_46_71), .A4(n_46_72), 
      .ZN(n_619));
   NAND2_X1 i_46_92 (.A1(n_599), .A2(multiplicand[19]), .ZN(n_46_73));
   NAND2_X1 i_46_93 (.A1(n_597), .A2(n_66), .ZN(n_46_74));
   NAND2_X1 i_46_94 (.A1(n_598), .A2(n_65), .ZN(n_46_75));
   NAND2_X1 i_46_95 (.A1(n_600), .A2(multiplicand[18]), .ZN(n_46_76));
   NAND4_X1 i_46_96 (.A1(n_46_73), .A2(n_46_74), .A3(n_46_75), .A4(n_46_76), 
      .ZN(n_620));
   NAND2_X1 i_46_97 (.A1(n_599), .A2(multiplicand[20]), .ZN(n_46_77));
   NAND2_X1 i_46_98 (.A1(n_597), .A2(n_67), .ZN(n_46_78));
   NAND2_X1 i_46_99 (.A1(n_598), .A2(n_66), .ZN(n_46_79));
   NAND2_X1 i_46_100 (.A1(n_600), .A2(multiplicand[19]), .ZN(n_46_80));
   NAND4_X1 i_46_101 (.A1(n_46_77), .A2(n_46_78), .A3(n_46_79), .A4(n_46_80), 
      .ZN(n_621));
   NAND2_X1 i_46_102 (.A1(n_599), .A2(multiplicand[21]), .ZN(n_46_81));
   NAND2_X1 i_46_103 (.A1(n_597), .A2(n_68), .ZN(n_46_82));
   NAND2_X1 i_46_104 (.A1(n_598), .A2(n_67), .ZN(n_46_83));
   NAND2_X1 i_46_105 (.A1(n_600), .A2(multiplicand[20]), .ZN(n_46_84));
   NAND4_X1 i_46_106 (.A1(n_46_81), .A2(n_46_82), .A3(n_46_83), .A4(n_46_84), 
      .ZN(n_622));
   NAND2_X1 i_46_107 (.A1(n_599), .A2(multiplicand[22]), .ZN(n_46_85));
   NAND2_X1 i_46_108 (.A1(n_597), .A2(n_69), .ZN(n_46_86));
   NAND2_X1 i_46_109 (.A1(n_598), .A2(n_68), .ZN(n_46_87));
   NAND2_X1 i_46_110 (.A1(n_600), .A2(multiplicand[21]), .ZN(n_46_88));
   NAND4_X1 i_46_111 (.A1(n_46_85), .A2(n_46_86), .A3(n_46_87), .A4(n_46_88), 
      .ZN(n_623));
   NAND2_X1 i_46_112 (.A1(n_599), .A2(multiplicand[23]), .ZN(n_46_89));
   NAND2_X1 i_46_113 (.A1(n_597), .A2(n_70), .ZN(n_46_90));
   NAND2_X1 i_46_114 (.A1(n_598), .A2(n_69), .ZN(n_46_91));
   NAND2_X1 i_46_115 (.A1(n_600), .A2(multiplicand[22]), .ZN(n_46_92));
   NAND4_X1 i_46_116 (.A1(n_46_89), .A2(n_46_90), .A3(n_46_91), .A4(n_46_92), 
      .ZN(n_624));
   NAND2_X1 i_46_117 (.A1(n_599), .A2(multiplicand[24]), .ZN(n_46_93));
   NAND2_X1 i_46_118 (.A1(n_597), .A2(n_71), .ZN(n_46_94));
   NAND2_X1 i_46_119 (.A1(n_598), .A2(n_70), .ZN(n_46_95));
   NAND2_X1 i_46_120 (.A1(n_600), .A2(multiplicand[23]), .ZN(n_46_96));
   NAND4_X1 i_46_121 (.A1(n_46_93), .A2(n_46_94), .A3(n_46_95), .A4(n_46_96), 
      .ZN(n_625));
   NAND2_X1 i_46_122 (.A1(n_599), .A2(multiplicand[25]), .ZN(n_46_97));
   NAND2_X1 i_46_123 (.A1(n_597), .A2(n_72), .ZN(n_46_98));
   NAND2_X1 i_46_124 (.A1(n_598), .A2(n_71), .ZN(n_46_99));
   NAND2_X1 i_46_125 (.A1(n_600), .A2(multiplicand[24]), .ZN(n_46_100));
   NAND4_X1 i_46_126 (.A1(n_46_97), .A2(n_46_98), .A3(n_46_99), .A4(n_46_100), 
      .ZN(n_626));
   NAND2_X1 i_46_127 (.A1(n_599), .A2(multiplicand[26]), .ZN(n_46_101));
   NAND2_X1 i_46_128 (.A1(n_597), .A2(n_73), .ZN(n_46_102));
   NAND2_X1 i_46_129 (.A1(n_598), .A2(n_72), .ZN(n_46_103));
   NAND2_X1 i_46_130 (.A1(n_600), .A2(multiplicand[25]), .ZN(n_46_104));
   NAND4_X1 i_46_131 (.A1(n_46_101), .A2(n_46_102), .A3(n_46_103), .A4(n_46_104), 
      .ZN(n_627));
   NAND2_X1 i_46_132 (.A1(n_599), .A2(multiplicand[27]), .ZN(n_46_105));
   NAND2_X1 i_46_133 (.A1(n_597), .A2(n_74), .ZN(n_46_106));
   NAND2_X1 i_46_134 (.A1(n_598), .A2(n_73), .ZN(n_46_107));
   NAND2_X1 i_46_135 (.A1(n_600), .A2(multiplicand[26]), .ZN(n_46_108));
   NAND4_X1 i_46_136 (.A1(n_46_105), .A2(n_46_106), .A3(n_46_107), .A4(n_46_108), 
      .ZN(n_628));
   NAND2_X1 i_46_137 (.A1(n_599), .A2(multiplicand[28]), .ZN(n_46_109));
   NAND2_X1 i_46_138 (.A1(n_597), .A2(n_75), .ZN(n_46_110));
   NAND2_X1 i_46_139 (.A1(n_598), .A2(n_74), .ZN(n_46_111));
   NAND2_X1 i_46_140 (.A1(n_600), .A2(multiplicand[27]), .ZN(n_46_112));
   NAND4_X1 i_46_141 (.A1(n_46_109), .A2(n_46_110), .A3(n_46_111), .A4(n_46_112), 
      .ZN(n_629));
   NAND2_X1 i_46_142 (.A1(n_599), .A2(multiplicand[29]), .ZN(n_46_113));
   NAND2_X1 i_46_143 (.A1(n_597), .A2(n_76), .ZN(n_46_114));
   NAND2_X1 i_46_144 (.A1(n_598), .A2(n_75), .ZN(n_46_115));
   NAND2_X1 i_46_145 (.A1(n_600), .A2(multiplicand[28]), .ZN(n_46_116));
   NAND4_X1 i_46_146 (.A1(n_46_113), .A2(n_46_114), .A3(n_46_115), .A4(n_46_116), 
      .ZN(n_630));
   NAND2_X1 i_46_147 (.A1(n_599), .A2(multiplicand[30]), .ZN(n_46_117));
   NAND2_X1 i_46_148 (.A1(n_597), .A2(n_77), .ZN(n_46_118));
   NAND2_X1 i_46_149 (.A1(n_598), .A2(n_76), .ZN(n_46_119));
   NAND2_X1 i_46_150 (.A1(n_600), .A2(multiplicand[29]), .ZN(n_46_120));
   NAND4_X1 i_46_151 (.A1(n_46_117), .A2(n_46_118), .A3(n_46_119), .A4(n_46_120), 
      .ZN(n_631));
   NAND2_X1 i_46_152 (.A1(n_599), .A2(multiplicand[31]), .ZN(n_46_121));
   NAND2_X1 i_46_153 (.A1(n_597), .A2(n_78), .ZN(n_46_122));
   NAND2_X1 i_46_154 (.A1(n_598), .A2(n_77), .ZN(n_46_123));
   NAND2_X1 i_46_155 (.A1(n_600), .A2(multiplicand[30]), .ZN(n_46_124));
   NAND4_X1 i_46_156 (.A1(n_46_121), .A2(n_46_122), .A3(n_46_123), .A4(n_46_124), 
      .ZN(n_632));
   NAND2_X1 i_46_157 (.A1(n_598), .A2(n_78), .ZN(n_46_125));
   NAND2_X1 i_46_158 (.A1(n_600), .A2(multiplicand[31]), .ZN(n_46_126));
   NAND4_X1 i_46_159 (.A1(n_46_121), .A2(n_46_122), .A3(n_46_125), .A4(n_46_126), 
      .ZN(n_633));
   INV_X1 i_47_0 (.A(n_45), .ZN(n_47_0));
   AND3_X1 i_47_1 (.A1(n_47_0), .A2(n_46), .A3(n_47), .ZN(n_634));
   INV_X1 i_47_2 (.A(n_47), .ZN(n_47_1));
   NOR3_X1 i_47_3 (.A1(n_47_1), .A2(n_47_0), .A3(n_46), .ZN(n_635));
   NOR3_X1 i_47_4 (.A1(n_47_0), .A2(n_46), .A3(n_47), .ZN(n_636));
   AOI22_X1 i_48_0 (.A1(multiplicand[0]), .A2(n_636), .B1(multiplicand[0]), 
      .B2(n_635), .ZN(n_48_0));
   INV_X1 i_48_1 (.A(n_48_0), .ZN(product[0]));
   AOI222_X1 i_48_2 (.A1(n_636), .A2(multiplicand[1]), .B1(n_635), .B2(n_48), 
      .C1(n_634), .C2(multiplicand[0]), .ZN(n_48_1));
   INV_X1 i_48_3 (.A(n_48_1), .ZN(product[1]));
   AOI222_X1 i_48_4 (.A1(n_636), .A2(multiplicand[2]), .B1(n_635), .B2(n_49), 
      .C1(n_634), .C2(n_48), .ZN(n_48_2));
   INV_X1 i_48_5 (.A(n_48_2), .ZN(n_637));
   AOI222_X1 i_48_6 (.A1(n_636), .A2(multiplicand[3]), .B1(n_635), .B2(n_50), 
      .C1(n_634), .C2(n_49), .ZN(n_48_3));
   INV_X1 i_48_7 (.A(n_48_3), .ZN(n_638));
   AOI222_X1 i_48_8 (.A1(n_636), .A2(multiplicand[4]), .B1(n_635), .B2(n_51), 
      .C1(n_634), .C2(n_50), .ZN(n_48_4));
   INV_X1 i_48_9 (.A(n_48_4), .ZN(n_639));
   AOI222_X1 i_48_10 (.A1(n_636), .A2(multiplicand[5]), .B1(n_635), .B2(n_52), 
      .C1(n_634), .C2(n_51), .ZN(n_48_5));
   INV_X1 i_48_11 (.A(n_48_5), .ZN(n_640));
   AOI222_X1 i_48_12 (.A1(n_636), .A2(multiplicand[6]), .B1(n_635), .B2(n_53), 
      .C1(n_634), .C2(n_52), .ZN(n_48_6));
   INV_X1 i_48_13 (.A(n_48_6), .ZN(n_641));
   AOI222_X1 i_48_14 (.A1(n_636), .A2(multiplicand[7]), .B1(n_635), .B2(n_54), 
      .C1(n_634), .C2(n_53), .ZN(n_48_7));
   INV_X1 i_48_15 (.A(n_48_7), .ZN(n_642));
   AOI222_X1 i_48_16 (.A1(n_636), .A2(multiplicand[8]), .B1(n_635), .B2(n_55), 
      .C1(n_634), .C2(n_54), .ZN(n_48_8));
   INV_X1 i_48_17 (.A(n_48_8), .ZN(n_643));
   AOI222_X1 i_48_18 (.A1(n_636), .A2(multiplicand[9]), .B1(n_635), .B2(n_56), 
      .C1(n_634), .C2(n_55), .ZN(n_48_9));
   INV_X1 i_48_19 (.A(n_48_9), .ZN(n_644));
   AOI222_X1 i_48_20 (.A1(n_636), .A2(multiplicand[10]), .B1(n_635), .B2(n_57), 
      .C1(n_634), .C2(n_56), .ZN(n_48_10));
   INV_X1 i_48_21 (.A(n_48_10), .ZN(n_645));
   AOI222_X1 i_48_22 (.A1(n_636), .A2(multiplicand[11]), .B1(n_635), .B2(n_58), 
      .C1(n_634), .C2(n_57), .ZN(n_48_11));
   INV_X1 i_48_23 (.A(n_48_11), .ZN(n_646));
   AOI222_X1 i_48_24 (.A1(n_636), .A2(multiplicand[12]), .B1(n_635), .B2(n_59), 
      .C1(n_634), .C2(n_58), .ZN(n_48_12));
   INV_X1 i_48_25 (.A(n_48_12), .ZN(n_647));
   AOI222_X1 i_48_26 (.A1(n_636), .A2(multiplicand[13]), .B1(n_635), .B2(n_60), 
      .C1(n_634), .C2(n_59), .ZN(n_48_13));
   INV_X1 i_48_27 (.A(n_48_13), .ZN(n_648));
   AOI222_X1 i_48_28 (.A1(n_636), .A2(multiplicand[14]), .B1(n_635), .B2(n_61), 
      .C1(n_634), .C2(n_60), .ZN(n_48_14));
   INV_X1 i_48_29 (.A(n_48_14), .ZN(n_649));
   AOI222_X1 i_48_30 (.A1(n_636), .A2(multiplicand[15]), .B1(n_635), .B2(n_62), 
      .C1(n_634), .C2(n_61), .ZN(n_48_15));
   INV_X1 i_48_31 (.A(n_48_15), .ZN(n_650));
   AOI222_X1 i_48_32 (.A1(n_636), .A2(multiplicand[16]), .B1(n_635), .B2(n_63), 
      .C1(n_634), .C2(n_62), .ZN(n_48_16));
   INV_X1 i_48_33 (.A(n_48_16), .ZN(n_651));
   AOI222_X1 i_48_34 (.A1(n_636), .A2(multiplicand[17]), .B1(n_635), .B2(n_64), 
      .C1(n_634), .C2(n_63), .ZN(n_48_17));
   INV_X1 i_48_35 (.A(n_48_17), .ZN(n_652));
   AOI222_X1 i_48_36 (.A1(n_636), .A2(multiplicand[18]), .B1(n_635), .B2(n_65), 
      .C1(n_634), .C2(n_64), .ZN(n_48_18));
   INV_X1 i_48_37 (.A(n_48_18), .ZN(n_653));
   AOI222_X1 i_48_38 (.A1(n_636), .A2(multiplicand[19]), .B1(n_635), .B2(n_66), 
      .C1(n_634), .C2(n_65), .ZN(n_48_19));
   INV_X1 i_48_39 (.A(n_48_19), .ZN(n_654));
   AOI222_X1 i_48_40 (.A1(n_636), .A2(multiplicand[20]), .B1(n_635), .B2(n_67), 
      .C1(n_634), .C2(n_66), .ZN(n_48_20));
   INV_X1 i_48_41 (.A(n_48_20), .ZN(n_655));
   AOI222_X1 i_48_42 (.A1(n_636), .A2(multiplicand[21]), .B1(n_635), .B2(n_68), 
      .C1(n_634), .C2(n_67), .ZN(n_48_21));
   INV_X1 i_48_43 (.A(n_48_21), .ZN(n_656));
   AOI222_X1 i_48_44 (.A1(n_636), .A2(multiplicand[22]), .B1(n_635), .B2(n_69), 
      .C1(n_634), .C2(n_68), .ZN(n_48_22));
   INV_X1 i_48_45 (.A(n_48_22), .ZN(n_657));
   AOI222_X1 i_48_46 (.A1(n_636), .A2(multiplicand[23]), .B1(n_635), .B2(n_70), 
      .C1(n_634), .C2(n_69), .ZN(n_48_23));
   INV_X1 i_48_47 (.A(n_48_23), .ZN(n_658));
   AOI222_X1 i_48_48 (.A1(n_636), .A2(multiplicand[24]), .B1(n_635), .B2(n_71), 
      .C1(n_634), .C2(n_70), .ZN(n_48_24));
   INV_X1 i_48_49 (.A(n_48_24), .ZN(n_659));
   AOI222_X1 i_48_50 (.A1(n_636), .A2(multiplicand[25]), .B1(n_635), .B2(n_72), 
      .C1(n_634), .C2(n_71), .ZN(n_48_25));
   INV_X1 i_48_51 (.A(n_48_25), .ZN(n_660));
   AOI222_X1 i_48_52 (.A1(n_636), .A2(multiplicand[26]), .B1(n_635), .B2(n_73), 
      .C1(n_634), .C2(n_72), .ZN(n_48_26));
   INV_X1 i_48_53 (.A(n_48_26), .ZN(n_661));
   AOI222_X1 i_48_54 (.A1(n_636), .A2(multiplicand[27]), .B1(n_635), .B2(n_74), 
      .C1(n_634), .C2(n_73), .ZN(n_48_27));
   INV_X1 i_48_55 (.A(n_48_27), .ZN(n_662));
   AOI222_X1 i_48_56 (.A1(n_636), .A2(multiplicand[28]), .B1(n_635), .B2(n_75), 
      .C1(n_634), .C2(n_74), .ZN(n_48_28));
   INV_X1 i_48_57 (.A(n_48_28), .ZN(n_663));
   AOI222_X1 i_48_58 (.A1(n_636), .A2(multiplicand[29]), .B1(n_635), .B2(n_76), 
      .C1(n_634), .C2(n_75), .ZN(n_48_29));
   INV_X1 i_48_59 (.A(n_48_29), .ZN(n_664));
   AOI222_X1 i_48_60 (.A1(n_636), .A2(multiplicand[30]), .B1(n_635), .B2(n_77), 
      .C1(n_634), .C2(n_76), .ZN(n_48_30));
   INV_X1 i_48_61 (.A(n_48_30), .ZN(n_665));
   NAND2_X1 i_48_62 (.A1(n_636), .A2(multiplicand[31]), .ZN(n_48_31));
   NAND2_X1 i_48_63 (.A1(n_635), .A2(n_78), .ZN(n_48_32));
   NAND2_X1 i_48_64 (.A1(n_634), .A2(n_77), .ZN(n_48_33));
   NAND3_X1 i_48_65 (.A1(n_48_31), .A2(n_48_32), .A3(n_48_33), .ZN(n_666));
   NAND2_X1 i_48_66 (.A1(n_634), .A2(n_78), .ZN(n_48_34));
   NAND3_X1 i_48_67 (.A1(n_48_31), .A2(n_48_32), .A3(n_48_34), .ZN(n_667));
   datapath__0_109 i_49 (.subRes({uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, 
      n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, n_106, 
      n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, n_97, n_96, n_95, 
      n_94, n_93, n_92, n_91, n_90, n_89, n_88, n_87, n_86, n_85, n_84, n_83, 
      1'b0, 1'b0}), .subRes0({uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, 
      uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, 
      uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, 
      n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, 
      n_142, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
      n_132, n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, 
      n_122, n_121, n_120, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes1({uc_57, uc_58, 
      uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, 
      uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, 
      uc_79, uc_80, uc_81, n_189, n_188, n_187, n_186, n_185, n_184, n_183, 
      n_182, n_181, n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, 
      n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
      n_162, n_161, n_160, n_159, n_158, n_157, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0}), .subRes2({uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, 
      uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, 
      uc_100, uc_101, uc_102, uc_103, uc_104, n_226, n_225, n_224, n_223, n_222, 
      n_221, n_220, n_219, n_218, n_217, n_216, n_215, n_214, n_213, n_212, 
      n_211, n_210, n_209, n_208, n_207, n_206, n_205, n_204, n_203, n_202, 
      n_201, n_200, n_199, n_198, n_197, n_196, n_195, n_194, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes3({uc_105, uc_106, uc_107, uc_108, 
      uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, 
      uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, n_263, 
      n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, n_253, 
      n_252, n_251, n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, 
      n_242, n_241, n_240, n_239, n_238, n_237, n_236, n_235, n_234, n_233, 
      n_232, n_231, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .subRes4({uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, 
      uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, 
      uc_143, uc_144, n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, 
      n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, n_284, n_283, 
      n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, 
      n_272, n_271, n_270, n_269, n_268, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes5({uc_145, uc_146, uc_147, 
      uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, uc_156, 
      uc_157, uc_158, uc_159, uc_160, uc_161, n_337, n_336, n_335, n_334, n_333, 
      n_332, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, n_323, 
      n_322, n_321, n_320, n_319, n_318, n_317, n_316, n_315, n_314, n_313, 
      n_312, n_311, n_310, n_309, n_308, n_307, n_306, n_305, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .subRes6({uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, 
      uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, n_374, n_373, 
      n_372, n_371, n_370, n_369, n_368, n_367, n_366, n_365, n_364, n_363, 
      n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, 
      n_352, n_351, n_350, n_349, n_348, n_347, n_346, n_345, n_344, n_343, 
      n_342, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes7({uc_177, uc_178, uc_179, uc_180, 
      uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, uc_189, 
      n_411, n_410, n_409, n_408, n_407, n_406, n_405, n_404, n_403, n_402, 
      n_401, n_400, n_399, n_398, n_397, n_396, n_395, n_394, n_393, n_392, 
      n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, n_383, n_382, 
      n_381, n_380, n_379, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes8({uc_190, 
      uc_191, uc_192, uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, 
      uc_200, n_448, n_447, n_446, n_445, n_444, n_443, n_442, n_441, n_440, 
      n_439, n_438, n_437, n_436, n_435, n_434, n_433, n_432, n_431, n_430, 
      n_429, n_428, n_427, n_426, n_425, n_424, n_423, n_422, n_421, n_420, 
      n_419, n_418, n_417, n_416, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .subRes9({uc_201, uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, 
      uc_209, n_485, n_484, n_483, n_482, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, n_468, n_467, 
      n_466, n_465, n_464, n_463, n_462, n_461, n_460, n_459, n_458, n_457, 
      n_456, n_455, n_454, n_453, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0}), .subRes10({uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, 
      uc_216, n_522, n_521, n_520, n_519, n_518, n_517, n_516, n_515, n_514, 
      n_513, n_512, n_511, n_510, n_509, n_508, n_507, n_506, n_505, n_504, 
      n_503, n_502, n_501, n_500, n_499, n_498, n_497, n_496, n_495, n_494, 
      n_493, n_492, n_491, n_490, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0}), .subRes11({uc_217, uc_218, uc_219, uc_220, 
      uc_221, n_559, n_558, n_557, n_556, n_555, n_554, n_553, n_552, n_551, 
      n_550, n_549, n_548, n_547, n_546, n_545, n_544, n_543, n_542, n_541, 
      n_540, n_539, n_538, n_537, n_536, n_535, n_534, n_533, n_532, n_531, 
      n_530, n_529, n_528, n_527, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes12({uc_222, uc_223, uc_224, 
      n_596, n_595, n_594, n_593, n_592, n_591, n_590, n_589, n_588, n_587, 
      n_586, n_585, n_584, n_583, n_582, n_581, n_580, n_579, n_578, n_577, 
      n_576, n_575, n_574, n_573, n_572, n_571, n_570, n_569, n_568, n_567, 
      n_566, n_565, n_564, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes13({uc_225, n_633, 
      n_632, n_631, n_630, n_629, n_628, n_627, n_626, n_625, n_624, n_623, 
      n_622, n_621, n_620, n_619, n_618, n_617, n_616, n_615, n_614, n_613, 
      n_612, n_611, n_610, n_609, n_608, n_607, n_606, n_605, n_604, n_603, 
      n_602, n_601, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .subRes14({uc_226, 
      uc_227, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, 
      uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, 
      uc_245, uc_246, uc_247, uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, 
      uc_254, uc_255, uc_256, n_667, n_666, n_665, n_664, n_663, n_662, n_661, 
      n_660, n_659, n_658, n_657, n_656, n_655, n_654, n_653, n_652, n_651, 
      n_650, n_649, n_648, n_647, n_646, n_645, n_644, n_643, n_642, n_641, 
      n_640, n_639, n_638, n_637, uc_257, uc_258}), .product_reg({product[63], 
      product[62], product[61], product[60], product[59], product[58], 
      product[57], product[56], product[55], product[54], product[53], 
      product[52], product[51], product[50], product[49], product[48], 
      product[47], product[46], product[45], product[44], product[43], 
      product[42], product[41], product[40], product[39], product[38], 
      product[37], product[36], product[35], product[34], product[33], 
      product[32], product[31], product[30], product[29], product[28], 
      product[27], product[26], product[25], product[24], product[23], 
      product[22], product[21], product[20], product[19], product[18], 
      product[17], product[16], product[15], product[14], product[13], 
      product[12], product[11], product[10], product[9], product[8], product[7], 
      product[6], product[5], product[4], product[3], product[2], uc_259, uc_260}));
endmodule

module RadixboothMult(i_clk, i_rst, i_en, i_inputA, i_inputB, o_result);
   input i_clk;
   input i_rst;
   input i_en;
   input [31:0]i_inputA;
   input [31:0]i_inputB;
   output [63:0]o_result;

   wire [31:0]B_reg;
   wire [31:0]A_reg;
   wire [63:0]out_reg;

   registerNbits_bbox_0 regB (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(
      i_inputB), .p_4(B_reg));
   registerNbits_bbox_1 outReg (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(
      out_reg), .p_4(o_result));
   registerNbits_bbox regA (.p_0(i_clk), .p_1(i_rst), .p_2(i_en), .p_3(i_inputA), 
      .p_4(A_reg));
   Radix4BoothMultiplier Radix4BoothMultiplierUnit (.multiplicand(A_reg), 
      .multiplier(B_reg), .product(out_reg));
endmodule
