module HA (
	input a,
	input b,
	output sum,
	output carry
);
assign {carry, sum} = a + b;
endmodule

module FA (
	input a,
	input b,
	input c,
	output sum,
	output carry
);
assign {carry, sum} = a + b + c;
endmodule

module signed_wallace_tree_multipler(
	input [31:0] A,
	input [31:0] B,
	output [63:0] result
);
reg [63:0] p[63:0];
// Set First 32 x 32 Products Of A x B
integer i;
always @(*) begin
	for(i = 0;i <= 63;i = i + 1)begin
		if(i >= 32)
			p[i] = {{32{B[31]}}, B} & {64{A[31]}};
		else
			p[i] = {{32{B[31]}}, B} & {64{A[i]}};
	end
end

wire [2232:0] r;
wire [2232:0] c;

HA HA_0(p[0][1], p[1][0], r[0], c[0]);
FA FA_0(p[0][2], p[1][1], p[2][0], r[1], c[1]);
FA FA_1(p[0][3], p[1][2], p[2][1], r[2], c[2]);
HA HA_1(p[3][0], c[1], r[3], c[3]);
FA FA_2(p[0][4], p[1][3], p[2][2], r[4], c[4]);
FA FA_3(p[0][5], p[1][4], p[2][3], r[5], c[5]);
FA FA_4(p[0][6], p[1][5], p[2][4], r[6], c[6]);
HA HA_2(p[3][3], p[4][2], r[7], c[7]);
FA FA_5(p[0][7], p[1][6], p[2][5], r[8], c[8]);
FA FA_6(p[0][8], p[1][7], p[2][6], r[9], c[9]);
FA FA_7(p[0][9], p[1][8], p[2][7], r[10], c[10]);
HA HA_3(p[3][6], p[4][5], r[11], c[11]);
FA FA_8(p[0][10], p[1][9], p[2][8], r[12], c[12]);
FA FA_9(p[3][7], p[4][6], p[5][5], r[13], c[13]);
FA FA_10(p[0][11], p[1][10], p[2][9], r[14], c[14]);
FA FA_11(p[3][8], p[4][7], p[5][6], r[15], c[15]);
HA HA_4(p[6][5], p[7][4], r[16], c[16]);
FA FA_12(p[0][12], p[1][11], p[2][10], r[17], c[17]);
FA FA_13(p[3][9], p[4][8], p[5][7], r[18], c[18]);
FA FA_14(p[0][13], p[1][12], p[2][11], r[19], c[19]);
FA FA_15(p[3][10], p[4][9], p[5][8], r[20], c[20]);
FA FA_16(p[0][14], p[1][13], p[2][12], r[21], c[21]);
FA FA_17(p[3][11], p[4][10], p[5][9], r[22], c[22]);
HA HA_5(p[6][8], p[7][7], r[23], c[23]);
FA FA_18(p[0][15], p[1][14], p[2][13], r[24], c[24]);
FA FA_19(p[3][12], p[4][11], p[5][10], r[25], c[25]);
FA FA_20(p[0][16], p[1][15], p[2][14], r[26], c[26]);
FA FA_21(p[3][13], p[4][12], p[5][11], r[27], c[27]);
FA FA_22(p[0][17], p[1][16], p[2][15], r[28], c[28]);
FA FA_23(p[3][14], p[4][13], p[5][12], r[29], c[29]);
HA HA_6(p[6][11], p[7][10], r[30], c[30]);
FA FA_24(p[0][18], p[1][17], p[2][16], r[31], c[31]);
FA FA_25(p[3][15], p[4][14], p[5][13], r[32], c[32]);
FA FA_26(p[6][12], p[7][11], p[8][10], r[33], c[33]);
FA FA_27(p[0][19], p[1][18], p[2][17], r[34], c[34]);
FA FA_28(p[3][16], p[4][15], p[5][14], r[35], c[35]);
FA FA_29(p[6][13], p[7][12], p[8][11], r[36], c[36]);
HA HA_7(p[9][10], p[10][9], r[37], c[37]);
FA FA_30(p[0][20], p[1][19], p[2][18], r[38], c[38]);
FA FA_31(p[3][17], p[4][16], p[5][15], r[39], c[39]);
FA FA_32(p[6][14], p[7][13], p[8][12], r[40], c[40]);
FA FA_33(p[0][21], p[1][20], p[2][19], r[41], c[41]);
FA FA_34(p[3][18], p[4][17], p[5][16], r[42], c[42]);
FA FA_35(p[6][15], p[7][14], p[8][13], r[43], c[43]);
FA FA_36(p[0][22], p[1][21], p[2][20], r[44], c[44]);
FA FA_37(p[3][19], p[4][18], p[5][17], r[45], c[45]);
FA FA_38(p[6][16], p[7][15], p[8][14], r[46], c[46]);
HA HA_8(p[9][13], p[10][12], r[47], c[47]);
FA FA_39(p[0][23], p[1][22], p[2][21], r[48], c[48]);
FA FA_40(p[3][20], p[4][19], p[5][18], r[49], c[49]);
FA FA_41(p[6][17], p[7][16], p[8][15], r[50], c[50]);
FA FA_42(p[0][24], p[1][23], p[2][22], r[51], c[51]);
FA FA_43(p[3][21], p[4][20], p[5][19], r[52], c[52]);
FA FA_44(p[6][18], p[7][17], p[8][16], r[53], c[53]);
FA FA_45(p[0][25], p[1][24], p[2][23], r[54], c[54]);
FA FA_46(p[3][22], p[4][21], p[5][20], r[55], c[55]);
FA FA_47(p[6][19], p[7][18], p[8][17], r[56], c[56]);
HA HA_9(p[9][16], p[10][15], r[57], c[57]);
FA FA_48(p[0][26], p[1][25], p[2][24], r[58], c[58]);
FA FA_49(p[3][23], p[4][22], p[5][21], r[59], c[59]);
FA FA_50(p[6][20], p[7][19], p[8][18], r[60], c[60]);
FA FA_51(p[9][17], p[10][16], p[11][15], r[61], c[61]);
FA FA_52(p[0][27], p[1][26], p[2][25], r[62], c[62]);
FA FA_53(p[3][24], p[4][23], p[5][22], r[63], c[63]);
FA FA_54(p[6][21], p[7][20], p[8][19], r[64], c[64]);
FA FA_55(p[9][18], p[10][17], p[11][16], r[65], c[65]);
HA HA_10(p[12][15], p[13][14], r[66], c[66]);
FA FA_56(p[0][28], p[1][27], p[2][26], r[67], c[67]);
FA FA_57(p[3][25], p[4][24], p[5][23], r[68], c[68]);
FA FA_58(p[6][22], p[7][21], p[8][20], r[69], c[69]);
FA FA_59(p[9][19], p[10][18], p[11][17], r[70], c[70]);
FA FA_60(p[0][29], p[1][28], p[2][27], r[71], c[71]);
FA FA_61(p[3][26], p[4][25], p[5][24], r[72], c[72]);
FA FA_62(p[6][23], p[7][22], p[8][21], r[73], c[73]);
FA FA_63(p[9][20], p[10][19], p[11][18], r[74], c[74]);
FA FA_64(p[0][30], p[1][29], p[2][28], r[75], c[75]);
FA FA_65(p[3][27], p[4][26], p[5][25], r[76], c[76]);
FA FA_66(p[6][24], p[7][23], p[8][22], r[77], c[77]);
FA FA_67(p[9][21], p[10][20], p[11][19], r[78], c[78]);
HA HA_11(p[12][18], p[13][17], r[79], c[79]);
FA FA_68(p[0][31], p[1][30], p[2][29], r[80], c[80]);
FA FA_69(p[3][28], p[4][27], p[5][26], r[81], c[81]);
FA FA_70(p[6][25], p[7][24], p[8][23], r[82], c[82]);
FA FA_71(p[9][22], p[10][21], p[11][20], r[83], c[83]);
FA FA_72(p[0][32], p[1][31], p[2][30], r[84], c[84]);
FA FA_73(p[3][29], p[4][28], p[5][27], r[85], c[85]);
FA FA_74(p[6][26], p[7][25], p[8][24], r[86], c[86]);
FA FA_75(p[9][23], p[10][22], p[11][21], r[87], c[87]);
FA FA_76(p[0][33], p[1][32], p[2][31], r[88], c[88]);
FA FA_77(p[3][30], p[4][29], p[5][28], r[89], c[89]);
FA FA_78(p[6][27], p[7][26], p[8][25], r[90], c[90]);
FA FA_79(p[9][24], p[10][23], p[11][22], r[91], c[91]);
HA HA_12(p[12][21], p[13][20], r[92], c[92]);
FA FA_80(p[0][34], p[1][33], p[2][32], r[93], c[93]);
FA FA_81(p[3][31], p[4][30], p[5][29], r[94], c[94]);
FA FA_82(p[6][28], p[7][27], p[8][26], r[95], c[95]);
FA FA_83(p[9][25], p[10][24], p[11][23], r[96], c[96]);
FA FA_84(p[12][22], p[13][21], p[14][20], r[97], c[97]);
FA FA_85(p[0][35], p[1][34], p[2][33], r[98], c[98]);
FA FA_86(p[3][32], p[4][31], p[5][30], r[99], c[99]);
FA FA_87(p[6][29], p[7][28], p[8][27], r[100], c[100]);
FA FA_88(p[9][26], p[10][25], p[11][24], r[101], c[101]);
FA FA_89(p[12][23], p[13][22], p[14][21], r[102], c[102]);
HA HA_13(p[15][20], p[16][19], r[103], c[103]);
FA FA_90(p[0][36], p[1][35], p[2][34], r[104], c[104]);
FA FA_91(p[3][33], p[4][32], p[5][31], r[105], c[105]);
FA FA_92(p[6][30], p[7][29], p[8][28], r[106], c[106]);
FA FA_93(p[9][27], p[10][26], p[11][25], r[107], c[107]);
FA FA_94(p[12][24], p[13][23], p[14][22], r[108], c[108]);
FA FA_95(p[0][37], p[1][36], p[2][35], r[109], c[109]);
FA FA_96(p[3][34], p[4][33], p[5][32], r[110], c[110]);
FA FA_97(p[6][31], p[7][30], p[8][29], r[111], c[111]);
FA FA_98(p[9][28], p[10][27], p[11][26], r[112], c[112]);
FA FA_99(p[12][25], p[13][24], p[14][23], r[113], c[113]);
FA FA_100(p[0][38], p[1][37], p[2][36], r[114], c[114]);
FA FA_101(p[3][35], p[4][34], p[5][33], r[115], c[115]);
FA FA_102(p[6][32], p[7][31], p[8][30], r[116], c[116]);
FA FA_103(p[9][29], p[10][28], p[11][27], r[117], c[117]);
FA FA_104(p[12][26], p[13][25], p[14][24], r[118], c[118]);
HA HA_14(p[15][23], p[16][22], r[119], c[119]);
FA FA_105(p[0][39], p[1][38], p[2][37], r[120], c[120]);
FA FA_106(p[3][36], p[4][35], p[5][34], r[121], c[121]);
FA FA_107(p[6][33], p[7][32], p[8][31], r[122], c[122]);
FA FA_108(p[9][30], p[10][29], p[11][28], r[123], c[123]);
FA FA_109(p[12][27], p[13][26], p[14][25], r[124], c[124]);
FA FA_110(p[0][40], p[1][39], p[2][38], r[125], c[125]);
FA FA_111(p[3][37], p[4][36], p[5][35], r[126], c[126]);
FA FA_112(p[6][34], p[7][33], p[8][32], r[127], c[127]);
FA FA_113(p[9][31], p[10][30], p[11][29], r[128], c[128]);
FA FA_114(p[12][28], p[13][27], p[14][26], r[129], c[129]);
FA FA_115(p[0][41], p[1][40], p[2][39], r[130], c[130]);
FA FA_116(p[3][38], p[4][37], p[5][36], r[131], c[131]);
FA FA_117(p[6][35], p[7][34], p[8][33], r[132], c[132]);
FA FA_118(p[9][32], p[10][31], p[11][30], r[133], c[133]);
FA FA_119(p[12][29], p[13][28], p[14][27], r[134], c[134]);
HA HA_15(p[15][26], p[16][25], r[135], c[135]);
FA FA_120(p[0][42], p[1][41], p[2][40], r[136], c[136]);
FA FA_121(p[3][39], p[4][38], p[5][37], r[137], c[137]);
FA FA_122(p[6][36], p[7][35], p[8][34], r[138], c[138]);
FA FA_123(p[9][33], p[10][32], p[11][31], r[139], c[139]);
FA FA_124(p[12][30], p[13][29], p[14][28], r[140], c[140]);
FA FA_125(p[15][27], p[16][26], p[17][25], r[141], c[141]);
FA FA_126(p[0][43], p[1][42], p[2][41], r[142], c[142]);
FA FA_127(p[3][40], p[4][39], p[5][38], r[143], c[143]);
FA FA_128(p[6][37], p[7][36], p[8][35], r[144], c[144]);
FA FA_129(p[9][34], p[10][33], p[11][32], r[145], c[145]);
FA FA_130(p[12][31], p[13][30], p[14][29], r[146], c[146]);
FA FA_131(p[15][28], p[16][27], p[17][26], r[147], c[147]);
HA HA_16(p[18][25], p[19][24], r[148], c[148]);
FA FA_132(p[0][44], p[1][43], p[2][42], r[149], c[149]);
FA FA_133(p[3][41], p[4][40], p[5][39], r[150], c[150]);
FA FA_134(p[6][38], p[7][37], p[8][36], r[151], c[151]);
FA FA_135(p[9][35], p[10][34], p[11][33], r[152], c[152]);
FA FA_136(p[12][32], p[13][31], p[14][30], r[153], c[153]);
FA FA_137(p[15][29], p[16][28], p[17][27], r[154], c[154]);
FA FA_138(p[0][45], p[1][44], p[2][43], r[155], c[155]);
FA FA_139(p[3][42], p[4][41], p[5][40], r[156], c[156]);
FA FA_140(p[6][39], p[7][38], p[8][37], r[157], c[157]);
FA FA_141(p[9][36], p[10][35], p[11][34], r[158], c[158]);
FA FA_142(p[12][33], p[13][32], p[14][31], r[159], c[159]);
FA FA_143(p[15][30], p[16][29], p[17][28], r[160], c[160]);
FA FA_144(p[0][46], p[1][45], p[2][44], r[161], c[161]);
FA FA_145(p[3][43], p[4][42], p[5][41], r[162], c[162]);
FA FA_146(p[6][40], p[7][39], p[8][38], r[163], c[163]);
FA FA_147(p[9][37], p[10][36], p[11][35], r[164], c[164]);
FA FA_148(p[12][34], p[13][33], p[14][32], r[165], c[165]);
FA FA_149(p[15][31], p[16][30], p[17][29], r[166], c[166]);
HA HA_17(p[18][28], p[19][27], r[167], c[167]);
FA FA_150(p[0][47], p[1][46], p[2][45], r[168], c[168]);
FA FA_151(p[3][44], p[4][43], p[5][42], r[169], c[169]);
FA FA_152(p[6][41], p[7][40], p[8][39], r[170], c[170]);
FA FA_153(p[9][38], p[10][37], p[11][36], r[171], c[171]);
FA FA_154(p[12][35], p[13][34], p[14][33], r[172], c[172]);
FA FA_155(p[15][32], p[16][31], p[17][30], r[173], c[173]);
FA FA_156(p[0][48], p[1][47], p[2][46], r[174], c[174]);
FA FA_157(p[3][45], p[4][44], p[5][43], r[175], c[175]);
FA FA_158(p[6][42], p[7][41], p[8][40], r[176], c[176]);
FA FA_159(p[9][39], p[10][38], p[11][37], r[177], c[177]);
FA FA_160(p[12][36], p[13][35], p[14][34], r[178], c[178]);
FA FA_161(p[15][33], p[16][32], p[17][31], r[179], c[179]);
FA FA_162(p[0][49], p[1][48], p[2][47], r[180], c[180]);
FA FA_163(p[3][46], p[4][45], p[5][44], r[181], c[181]);
FA FA_164(p[6][43], p[7][42], p[8][41], r[182], c[182]);
FA FA_165(p[9][40], p[10][39], p[11][38], r[183], c[183]);
FA FA_166(p[12][37], p[13][36], p[14][35], r[184], c[184]);
FA FA_167(p[15][34], p[16][33], p[17][32], r[185], c[185]);
HA HA_18(p[18][31], p[19][30], r[186], c[186]);
FA FA_168(p[0][50], p[1][49], p[2][48], r[187], c[187]);
FA FA_169(p[3][47], p[4][46], p[5][45], r[188], c[188]);
FA FA_170(p[6][44], p[7][43], p[8][42], r[189], c[189]);
FA FA_171(p[9][41], p[10][40], p[11][39], r[190], c[190]);
FA FA_172(p[12][38], p[13][37], p[14][36], r[191], c[191]);
FA FA_173(p[15][35], p[16][34], p[17][33], r[192], c[192]);
FA FA_174(p[18][32], p[19][31], p[20][30], r[193], c[193]);
FA FA_175(p[0][51], p[1][50], p[2][49], r[194], c[194]);
FA FA_176(p[3][48], p[4][47], p[5][46], r[195], c[195]);
FA FA_177(p[6][45], p[7][44], p[8][43], r[196], c[196]);
FA FA_178(p[9][42], p[10][41], p[11][40], r[197], c[197]);
FA FA_179(p[12][39], p[13][38], p[14][37], r[198], c[198]);
FA FA_180(p[15][36], p[16][35], p[17][34], r[199], c[199]);
FA FA_181(p[18][33], p[19][32], p[20][31], r[200], c[200]);
HA HA_19(p[21][30], p[22][29], r[201], c[201]);
FA FA_182(p[0][52], p[1][51], p[2][50], r[202], c[202]);
FA FA_183(p[3][49], p[4][48], p[5][47], r[203], c[203]);
FA FA_184(p[6][46], p[7][45], p[8][44], r[204], c[204]);
FA FA_185(p[9][43], p[10][42], p[11][41], r[205], c[205]);
FA FA_186(p[12][40], p[13][39], p[14][38], r[206], c[206]);
FA FA_187(p[15][37], p[16][36], p[17][35], r[207], c[207]);
FA FA_188(p[18][34], p[19][33], p[20][32], r[208], c[208]);
FA FA_189(p[0][53], p[1][52], p[2][51], r[209], c[209]);
FA FA_190(p[3][50], p[4][49], p[5][48], r[210], c[210]);
FA FA_191(p[6][47], p[7][46], p[8][45], r[211], c[211]);
FA FA_192(p[9][44], p[10][43], p[11][42], r[212], c[212]);
FA FA_193(p[12][41], p[13][40], p[14][39], r[213], c[213]);
FA FA_194(p[15][38], p[16][37], p[17][36], r[214], c[214]);
FA FA_195(p[18][35], p[19][34], p[20][33], r[215], c[215]);
FA FA_196(p[0][54], p[1][53], p[2][52], r[216], c[216]);
FA FA_197(p[3][51], p[4][50], p[5][49], r[217], c[217]);
FA FA_198(p[6][48], p[7][47], p[8][46], r[218], c[218]);
FA FA_199(p[9][45], p[10][44], p[11][43], r[219], c[219]);
FA FA_200(p[12][42], p[13][41], p[14][40], r[220], c[220]);
FA FA_201(p[15][39], p[16][38], p[17][37], r[221], c[221]);
FA FA_202(p[18][36], p[19][35], p[20][34], r[222], c[222]);
HA HA_20(p[21][33], p[22][32], r[223], c[223]);
FA FA_203(p[0][55], p[1][54], p[2][53], r[224], c[224]);
FA FA_204(p[3][52], p[4][51], p[5][50], r[225], c[225]);
FA FA_205(p[6][49], p[7][48], p[8][47], r[226], c[226]);
FA FA_206(p[9][46], p[10][45], p[11][44], r[227], c[227]);
FA FA_207(p[12][43], p[13][42], p[14][41], r[228], c[228]);
FA FA_208(p[15][40], p[16][39], p[17][38], r[229], c[229]);
FA FA_209(p[18][37], p[19][36], p[20][35], r[230], c[230]);
FA FA_210(p[0][56], p[1][55], p[2][54], r[231], c[231]);
FA FA_211(p[3][53], p[4][52], p[5][51], r[232], c[232]);
FA FA_212(p[6][50], p[7][49], p[8][48], r[233], c[233]);
FA FA_213(p[9][47], p[10][46], p[11][45], r[234], c[234]);
FA FA_214(p[12][44], p[13][43], p[14][42], r[235], c[235]);
FA FA_215(p[15][41], p[16][40], p[17][39], r[236], c[236]);
FA FA_216(p[18][38], p[19][37], p[20][36], r[237], c[237]);
FA FA_217(p[0][57], p[1][56], p[2][55], r[238], c[238]);
FA FA_218(p[3][54], p[4][53], p[5][52], r[239], c[239]);
FA FA_219(p[6][51], p[7][50], p[8][49], r[240], c[240]);
FA FA_220(p[9][48], p[10][47], p[11][46], r[241], c[241]);
FA FA_221(p[12][45], p[13][44], p[14][43], r[242], c[242]);
FA FA_222(p[15][42], p[16][41], p[17][40], r[243], c[243]);
FA FA_223(p[18][39], p[19][38], p[20][37], r[244], c[244]);
HA HA_21(p[21][36], p[22][35], r[245], c[245]);
FA FA_224(p[0][58], p[1][57], p[2][56], r[246], c[246]);
FA FA_225(p[3][55], p[4][54], p[5][53], r[247], c[247]);
FA FA_226(p[6][52], p[7][51], p[8][50], r[248], c[248]);
FA FA_227(p[9][49], p[10][48], p[11][47], r[249], c[249]);
FA FA_228(p[12][46], p[13][45], p[14][44], r[250], c[250]);
FA FA_229(p[15][43], p[16][42], p[17][41], r[251], c[251]);
FA FA_230(p[18][40], p[19][39], p[20][38], r[252], c[252]);
FA FA_231(p[21][37], p[22][36], p[23][35], r[253], c[253]);
FA FA_232(p[0][59], p[1][58], p[2][57], r[254], c[254]);
FA FA_233(p[3][56], p[4][55], p[5][54], r[255], c[255]);
FA FA_234(p[6][53], p[7][52], p[8][51], r[256], c[256]);
FA FA_235(p[9][50], p[10][49], p[11][48], r[257], c[257]);
FA FA_236(p[12][47], p[13][46], p[14][45], r[258], c[258]);
FA FA_237(p[15][44], p[16][43], p[17][42], r[259], c[259]);
FA FA_238(p[18][41], p[19][40], p[20][39], r[260], c[260]);
FA FA_239(p[21][38], p[22][37], p[23][36], r[261], c[261]);
HA HA_22(p[24][35], p[25][34], r[262], c[262]);
FA FA_240(p[0][60], p[1][59], p[2][58], r[263], c[263]);
FA FA_241(p[3][57], p[4][56], p[5][55], r[264], c[264]);
FA FA_242(p[6][54], p[7][53], p[8][52], r[265], c[265]);
FA FA_243(p[9][51], p[10][50], p[11][49], r[266], c[266]);
FA FA_244(p[12][48], p[13][47], p[14][46], r[267], c[267]);
FA FA_245(p[15][45], p[16][44], p[17][43], r[268], c[268]);
FA FA_246(p[18][42], p[19][41], p[20][40], r[269], c[269]);
FA FA_247(p[21][39], p[22][38], p[23][37], r[270], c[270]);
FA FA_248(p[0][61], p[1][60], p[2][59], r[271], c[271]);
FA FA_249(p[3][58], p[4][57], p[5][56], r[272], c[272]);
FA FA_250(p[6][55], p[7][54], p[8][53], r[273], c[273]);
FA FA_251(p[9][52], p[10][51], p[11][50], r[274], c[274]);
FA FA_252(p[12][49], p[13][48], p[14][47], r[275], c[275]);
FA FA_253(p[15][46], p[16][45], p[17][44], r[276], c[276]);
FA FA_254(p[18][43], p[19][42], p[20][41], r[277], c[277]);
FA FA_255(p[21][40], p[22][39], p[23][38], r[278], c[278]);
FA FA_256(p[0][62], p[1][61], p[2][60], r[279], c[279]);
FA FA_257(p[3][59], p[4][58], p[5][57], r[280], c[280]);
FA FA_258(p[6][56], p[7][55], p[8][54], r[281], c[281]);
FA FA_259(p[9][53], p[10][52], p[11][51], r[282], c[282]);
FA FA_260(p[12][50], p[13][49], p[14][48], r[283], c[283]);
FA FA_261(p[15][47], p[16][46], p[17][45], r[284], c[284]);
FA FA_262(p[18][44], p[19][43], p[20][42], r[285], c[285]);
FA FA_263(p[21][41], p[22][40], p[23][39], r[286], c[286]);
HA HA_23(p[24][38], p[25][37], r[287], c[287]);
FA FA_264(p[0][63], p[1][62], p[2][61], r[288], c[288]);
FA FA_265(p[3][60], p[4][59], p[5][58], r[289], c[289]);
FA FA_266(p[6][57], p[7][56], p[8][55], r[290], c[290]);
FA FA_267(p[9][54], p[10][53], p[11][52], r[291], c[291]);
FA FA_268(p[12][51], p[13][50], p[14][49], r[292], c[292]);
FA FA_269(p[15][48], p[16][47], p[17][46], r[293], c[293]);
FA FA_270(p[18][45], p[19][44], p[20][43], r[294], c[294]);
FA FA_271(p[21][42], p[22][41], p[23][40], r[295], c[295]);
HA HA_24(c[0], r[1], r[296], c[296]);
FA FA_272(r[2], r[3], c[296], r[297], c[297]);
FA FA_273(p[3][1], p[4][0], c[2], r[298], c[298]);
FA FA_274(p[3][2], p[4][1], p[5][0], r[299], c[299]);
FA FA_275(p[5][1], p[6][0], c[5], r[300], c[300]);
FA FA_276(p[3][4], p[4][3], p[5][2], r[301], c[301]);
FA FA_277(p[3][5], p[4][4], p[5][3], r[302], c[302]);
FA FA_278(p[5][4], p[6][3], p[7][2], r[303], c[303]);
FA FA_279(p[6][4], p[7][3], p[8][2], r[304], c[304]);
FA FA_280(p[8][3], p[9][2], p[10][1], r[305], c[305]);
FA FA_281(p[6][6], p[7][5], p[8][4], r[306], c[306]);
FA FA_282(p[9][3], p[10][2], p[11][1], r[307], c[307]);
FA FA_283(p[6][7], p[7][6], p[8][5], r[308], c[308]);
FA FA_284(p[9][4], p[10][3], p[11][2], r[309], c[309]);
HA HA_25(p[12][1], p[13][0], r[310], c[310]);
FA FA_285(p[8][6], p[9][5], p[10][4], r[311], c[311]);
FA FA_286(p[11][3], p[12][2], p[13][1], r[312], c[312]);
FA FA_287(p[6][9], p[7][8], p[8][7], r[313], c[313]);
FA FA_288(p[9][6], p[10][5], p[11][4], r[314], c[314]);
HA HA_26(p[12][3], p[13][2], r[315], c[315]);
FA FA_289(p[6][10], p[7][9], p[8][8], r[316], c[316]);
FA FA_290(p[9][7], p[10][6], p[11][5], r[317], c[317]);
FA FA_291(p[8][9], p[9][8], p[10][7], r[318], c[318]);
FA FA_292(p[11][6], p[12][5], p[13][4], r[319], c[319]);
HA HA_27(p[14][3], p[15][2], r[320], c[320]);
FA FA_293(p[9][9], p[10][8], p[11][7], r[321], c[321]);
FA FA_294(p[12][6], p[13][5], p[14][4], r[322], c[322]);
FA FA_295(p[11][8], p[12][7], p[13][6], r[323], c[323]);
FA FA_296(p[14][5], p[15][4], p[16][3], r[324], c[324]);
FA FA_297(p[9][11], p[10][10], p[11][9], r[325], c[325]);
FA FA_298(p[12][8], p[13][7], p[14][6], r[326], c[326]);
FA FA_299(p[15][5], p[16][4], p[17][3], r[327], c[327]);
FA FA_300(p[9][12], p[10][11], p[11][10], r[328], c[328]);
FA FA_301(p[12][9], p[13][8], p[14][7], r[329], c[329]);
FA FA_302(p[15][6], p[16][5], p[17][4], r[330], c[330]);
FA FA_303(p[11][11], p[12][10], p[13][9], r[331], c[331]);
FA FA_304(p[14][8], p[15][7], p[16][6], r[332], c[332]);
FA FA_305(p[17][5], p[18][4], p[19][3], r[333], c[333]);
FA FA_306(p[9][14], p[10][13], p[11][12], r[334], c[334]);
FA FA_307(p[12][11], p[13][10], p[14][9], r[335], c[335]);
FA FA_308(p[15][8], p[16][7], p[17][6], r[336], c[336]);
FA FA_309(p[9][15], p[10][14], p[11][13], r[337], c[337]);
FA FA_310(p[12][12], p[13][11], p[14][10], r[338], c[338]);
FA FA_311(p[15][9], p[16][8], p[17][7], r[339], c[339]);
FA FA_312(p[11][14], p[12][13], p[13][12], r[340], c[340]);
FA FA_313(p[14][11], p[15][10], p[16][9], r[341], c[341]);
FA FA_314(p[17][8], p[18][7], p[19][6], r[342], c[342]);
FA FA_315(p[12][14], p[13][13], p[14][12], r[343], c[343]);
FA FA_316(p[15][11], p[16][10], p[17][9], r[344], c[344]);
FA FA_317(p[18][8], p[19][7], p[20][6], r[345], c[345]);
HA HA_28(p[21][5], p[22][4], r[346], c[346]);
FA FA_318(p[14][13], p[15][12], p[16][11], r[347], c[347]);
FA FA_319(p[17][10], p[18][9], p[19][8], r[348], c[348]);
FA FA_320(p[20][7], p[21][6], p[22][5], r[349], c[349]);
FA FA_321(p[12][16], p[13][15], p[14][14], r[350], c[350]);
FA FA_322(p[15][13], p[16][12], p[17][11], r[351], c[351]);
FA FA_323(p[18][10], p[19][9], p[20][8], r[352], c[352]);
HA HA_29(p[21][7], p[22][6], r[353], c[353]);
FA FA_324(p[12][17], p[13][16], p[14][15], r[354], c[354]);
FA FA_325(p[15][14], p[16][13], p[17][12], r[355], c[355]);
FA FA_326(p[18][11], p[19][10], p[20][9], r[356], c[356]);
FA FA_327(p[21][8], p[22][7], p[23][6], r[357], c[357]);
FA FA_328(p[14][16], p[15][15], p[16][14], r[358], c[358]);
FA FA_329(p[17][13], p[18][12], p[19][11], r[359], c[359]);
FA FA_330(p[20][10], p[21][9], p[22][8], r[360], c[360]);
FA FA_331(p[23][7], p[24][6], p[25][5], r[361], c[361]);
FA FA_332(p[12][19], p[13][18], p[14][17], r[362], c[362]);
FA FA_333(p[15][16], p[16][15], p[17][14], r[363], c[363]);
FA FA_334(p[18][13], p[19][12], p[20][11], r[364], c[364]);
FA FA_335(p[21][10], p[22][9], p[23][8], r[365], c[365]);
FA FA_336(p[12][20], p[13][19], p[14][18], r[366], c[366]);
FA FA_337(p[15][17], p[16][16], p[17][15], r[367], c[367]);
FA FA_338(p[18][14], p[19][13], p[20][12], r[368], c[368]);
FA FA_339(p[21][11], p[22][10], p[23][9], r[369], c[369]);
FA FA_340(p[14][19], p[15][18], p[16][17], r[370], c[370]);
FA FA_341(p[17][16], p[18][15], p[19][14], r[371], c[371]);
FA FA_342(p[20][13], p[21][12], p[22][11], r[372], c[372]);
FA FA_343(p[23][10], p[24][9], p[25][8], r[373], c[373]);
FA FA_344(p[15][19], p[16][18], p[17][17], r[374], c[374]);
FA FA_345(p[18][16], p[19][15], p[20][14], r[375], c[375]);
FA FA_346(p[21][13], p[22][12], p[23][11], r[376], c[376]);
FA FA_347(p[24][10], p[25][9], p[26][8], r[377], c[377]);
FA FA_348(p[17][18], p[18][17], p[19][16], r[378], c[378]);
FA FA_349(p[20][15], p[21][14], p[22][13], r[379], c[379]);
FA FA_350(p[23][12], p[24][11], p[25][10], r[380], c[380]);
FA FA_351(p[26][9], p[27][8], p[28][7], r[381], c[381]);
FA FA_352(p[15][21], p[16][20], p[17][19], r[382], c[382]);
FA FA_353(p[18][18], p[19][17], p[20][16], r[383], c[383]);
FA FA_354(p[21][15], p[22][14], p[23][13], r[384], c[384]);
FA FA_355(p[24][12], p[25][11], p[26][10], r[385], c[385]);
FA FA_356(p[15][22], p[16][21], p[17][20], r[386], c[386]);
FA FA_357(p[18][19], p[19][18], p[20][17], r[387], c[387]);
FA FA_358(p[21][16], p[22][15], p[23][14], r[388], c[388]);
FA FA_359(p[24][13], p[25][12], p[26][11], r[389], c[389]);
FA FA_360(p[17][21], p[18][20], p[19][19], r[390], c[390]);
FA FA_361(p[20][18], p[21][17], p[22][16], r[391], c[391]);
FA FA_362(p[23][15], p[24][14], p[25][13], r[392], c[392]);
FA FA_363(p[26][12], p[27][11], p[28][10], r[393], c[393]);
FA FA_364(p[15][24], p[16][23], p[17][22], r[394], c[394]);
FA FA_365(p[18][21], p[19][20], p[20][19], r[395], c[395]);
FA FA_366(p[21][18], p[22][17], p[23][16], r[396], c[396]);
FA FA_367(p[24][15], p[25][14], p[26][13], r[397], c[397]);
FA FA_368(p[27][12], p[28][11], p[29][10], r[398], c[398]);
FA FA_369(p[15][25], p[16][24], p[17][23], r[399], c[399]);
FA FA_370(p[18][22], p[19][21], p[20][20], r[400], c[400]);
FA FA_371(p[21][19], p[22][18], p[23][17], r[401], c[401]);
FA FA_372(p[24][16], p[25][15], p[26][14], r[402], c[402]);
FA FA_373(p[27][13], p[28][12], p[29][11], r[403], c[403]);
HA HA_30(p[30][10], p[31][9], r[404], c[404]);
FA FA_374(p[17][24], p[18][23], p[19][22], r[405], c[405]);
FA FA_375(p[20][21], p[21][20], p[22][19], r[406], c[406]);
FA FA_376(p[23][18], p[24][17], p[25][16], r[407], c[407]);
FA FA_377(p[26][15], p[27][14], p[28][13], r[408], c[408]);
FA FA_378(p[29][12], p[30][11], p[31][10], r[409], c[409]);
FA FA_379(p[18][24], p[19][23], p[20][22], r[410], c[410]);
FA FA_380(p[21][21], p[22][20], p[23][19], r[411], c[411]);
FA FA_381(p[24][18], p[25][17], p[26][16], r[412], c[412]);
FA FA_382(p[27][15], p[28][14], p[29][13], r[413], c[413]);
FA FA_383(p[30][12], p[31][11], p[32][10], r[414], c[414]);
FA FA_384(p[20][23], p[21][22], p[22][21], r[415], c[415]);
FA FA_385(p[23][20], p[24][19], p[25][18], r[416], c[416]);
FA FA_386(p[26][17], p[27][16], p[28][15], r[417], c[417]);
FA FA_387(p[29][14], p[30][13], p[31][12], r[418], c[418]);
FA FA_388(p[32][11], p[33][10], p[34][9], r[419], c[419]);
FA FA_389(p[18][26], p[19][25], p[20][24], r[420], c[420]);
FA FA_390(p[21][23], p[22][22], p[23][21], r[421], c[421]);
FA FA_391(p[24][20], p[25][19], p[26][18], r[422], c[422]);
FA FA_392(p[27][17], p[28][16], p[29][15], r[423], c[423]);
FA FA_393(p[30][14], p[31][13], p[32][12], r[424], c[424]);
FA FA_394(p[18][27], p[19][26], p[20][25], r[425], c[425]);
FA FA_395(p[21][24], p[22][23], p[23][22], r[426], c[426]);
FA FA_396(p[24][21], p[25][20], p[26][19], r[427], c[427]);
FA FA_397(p[27][18], p[28][17], p[29][16], r[428], c[428]);
FA FA_398(p[30][15], p[31][14], p[32][13], r[429], c[429]);
FA FA_399(p[20][26], p[21][25], p[22][24], r[430], c[430]);
FA FA_400(p[23][23], p[24][22], p[25][21], r[431], c[431]);
FA FA_401(p[26][20], p[27][19], p[28][18], r[432], c[432]);
FA FA_402(p[29][17], p[30][16], p[31][15], r[433], c[433]);
FA FA_403(p[32][14], p[33][13], p[34][12], r[434], c[434]);
FA FA_404(p[18][29], p[19][28], p[20][27], r[435], c[435]);
FA FA_405(p[21][26], p[22][25], p[23][24], r[436], c[436]);
FA FA_406(p[24][23], p[25][22], p[26][21], r[437], c[437]);
FA FA_407(p[27][20], p[28][19], p[29][18], r[438], c[438]);
FA FA_408(p[30][17], p[31][16], p[32][15], r[439], c[439]);
FA FA_409(p[33][14], p[34][13], p[35][12], r[440], c[440]);
FA FA_410(p[18][30], p[19][29], p[20][28], r[441], c[441]);
FA FA_411(p[21][27], p[22][26], p[23][25], r[442], c[442]);
FA FA_412(p[24][24], p[25][23], p[26][22], r[443], c[443]);
FA FA_413(p[27][21], p[28][20], p[29][19], r[444], c[444]);
FA FA_414(p[30][18], p[31][17], p[32][16], r[445], c[445]);
FA FA_415(p[33][15], p[34][14], p[35][13], r[446], c[446]);
FA FA_416(p[20][29], p[21][28], p[22][27], r[447], c[447]);
FA FA_417(p[23][26], p[24][25], p[25][24], r[448], c[448]);
FA FA_418(p[26][23], p[27][22], p[28][21], r[449], c[449]);
FA FA_419(p[29][20], p[30][19], p[31][18], r[450], c[450]);
FA FA_420(p[32][17], p[33][16], p[34][15], r[451], c[451]);
FA FA_421(p[35][14], p[36][13], p[37][12], r[452], c[452]);
FA FA_422(p[21][29], p[22][28], p[23][27], r[453], c[453]);
FA FA_423(p[24][26], p[25][25], p[26][24], r[454], c[454]);
FA FA_424(p[27][23], p[28][22], p[29][21], r[455], c[455]);
FA FA_425(p[30][20], p[31][19], p[32][18], r[456], c[456]);
FA FA_426(p[33][17], p[34][16], p[35][15], r[457], c[457]);
FA FA_427(p[36][14], p[37][13], p[38][12], r[458], c[458]);
HA HA_31(p[39][11], p[40][10], r[459], c[459]);
FA FA_428(p[23][28], p[24][27], p[25][26], r[460], c[460]);
FA FA_429(p[26][25], p[27][24], p[28][23], r[461], c[461]);
FA FA_430(p[29][22], p[30][21], p[31][20], r[462], c[462]);
FA FA_431(p[32][19], p[33][18], p[34][17], r[463], c[463]);
FA FA_432(p[35][16], p[36][15], p[37][14], r[464], c[464]);
FA FA_433(p[38][13], p[39][12], p[40][11], r[465], c[465]);
FA FA_434(p[21][31], p[22][30], p[23][29], r[466], c[466]);
FA FA_435(p[24][28], p[25][27], p[26][26], r[467], c[467]);
FA FA_436(p[27][25], p[28][24], p[29][23], r[468], c[468]);
FA FA_437(p[30][22], p[31][21], p[32][20], r[469], c[469]);
FA FA_438(p[33][19], p[34][18], p[35][17], r[470], c[470]);
FA FA_439(p[36][16], p[37][15], p[38][14], r[471], c[471]);
HA HA_32(p[39][13], p[40][12], r[472], c[472]);
FA FA_440(p[21][32], p[22][31], p[23][30], r[473], c[473]);
FA FA_441(p[24][29], p[25][28], p[26][27], r[474], c[474]);
FA FA_442(p[27][26], p[28][25], p[29][24], r[475], c[475]);
FA FA_443(p[30][23], p[31][22], p[32][21], r[476], c[476]);
FA FA_444(p[33][20], p[34][19], p[35][18], r[477], c[477]);
FA FA_445(p[36][17], p[37][16], p[38][15], r[478], c[478]);
FA FA_446(p[23][31], p[24][30], p[25][29], r[479], c[479]);
FA FA_447(p[26][28], p[27][27], p[28][26], r[480], c[480]);
FA FA_448(p[29][25], p[30][24], p[31][23], r[481], c[481]);
FA FA_449(p[32][22], p[33][21], p[34][20], r[482], c[482]);
FA FA_450(p[35][19], p[36][18], p[37][17], r[483], c[483]);
FA FA_451(p[38][16], p[39][15], p[40][14], r[484], c[484]);
HA HA_33(p[41][13], p[42][12], r[485], c[485]);
FA FA_452(p[21][34], p[22][33], p[23][32], r[486], c[486]);
FA FA_453(p[24][31], p[25][30], p[26][29], r[487], c[487]);
FA FA_454(p[27][28], p[28][27], p[29][26], r[488], c[488]);
FA FA_455(p[30][25], p[31][24], p[32][23], r[489], c[489]);
FA FA_456(p[33][22], p[34][21], p[35][20], r[490], c[490]);
FA FA_457(p[36][19], p[37][18], p[38][17], r[491], c[491]);
FA FA_458(p[39][16], p[40][15], p[41][14], r[492], c[492]);
FA FA_459(p[21][35], p[22][34], p[23][33], r[493], c[493]);
FA FA_460(p[24][32], p[25][31], p[26][30], r[494], c[494]);
FA FA_461(p[27][29], p[28][28], p[29][27], r[495], c[495]);
FA FA_462(p[30][26], p[31][25], p[32][24], r[496], c[496]);
FA FA_463(p[33][23], p[34][22], p[35][21], r[497], c[497]);
FA FA_464(p[36][20], p[37][19], p[38][18], r[498], c[498]);
FA FA_465(p[39][17], p[40][16], p[41][15], r[499], c[499]);
FA FA_466(p[23][34], p[24][33], p[25][32], r[500], c[500]);
FA FA_467(p[26][31], p[27][30], p[28][29], r[501], c[501]);
FA FA_468(p[29][28], p[30][27], p[31][26], r[502], c[502]);
FA FA_469(p[32][25], p[33][24], p[34][23], r[503], c[503]);
FA FA_470(p[35][22], p[36][21], p[37][20], r[504], c[504]);
FA FA_471(p[38][19], p[39][18], p[40][17], r[505], c[505]);
FA FA_472(p[41][16], p[42][15], p[43][14], r[506], c[506]);
FA FA_473(p[24][34], p[25][33], p[26][32], r[507], c[507]);
FA FA_474(p[27][31], p[28][30], p[29][29], r[508], c[508]);
FA FA_475(p[30][28], p[31][27], p[32][26], r[509], c[509]);
FA FA_476(p[33][25], p[34][24], p[35][23], r[510], c[510]);
FA FA_477(p[36][22], p[37][21], p[38][20], r[511], c[511]);
FA FA_478(p[39][19], p[40][18], p[41][17], r[512], c[512]);
FA FA_479(p[42][16], p[43][15], p[44][14], r[513], c[513]);
FA FA_480(p[26][33], p[27][32], p[28][31], r[514], c[514]);
FA FA_481(p[29][30], p[30][29], p[31][28], r[515], c[515]);
FA FA_482(p[32][27], p[33][26], p[34][25], r[516], c[516]);
FA FA_483(p[35][24], p[36][23], p[37][22], r[517], c[517]);
FA FA_484(p[38][21], p[39][20], p[40][19], r[518], c[518]);
FA FA_485(p[41][18], p[42][17], p[43][16], r[519], c[519]);
FA FA_486(p[44][15], p[45][14], p[46][13], r[520], c[520]);
FA FA_487(p[24][36], p[25][35], p[26][34], r[521], c[521]);
FA FA_488(p[27][33], p[28][32], p[29][31], r[522], c[522]);
FA FA_489(p[30][30], p[31][29], p[32][28], r[523], c[523]);
FA FA_490(p[33][27], p[34][26], p[35][25], r[524], c[524]);
FA FA_491(p[36][24], p[37][23], p[38][22], r[525], c[525]);
FA FA_492(p[39][21], p[40][20], p[41][19], r[526], c[526]);
FA FA_493(p[42][18], p[43][17], p[44][16], r[527], c[527]);
FA FA_494(p[24][37], p[25][36], p[26][35], r[528], c[528]);
FA FA_495(p[27][34], p[28][33], p[29][32], r[529], c[529]);
FA FA_496(p[30][31], p[31][30], p[32][29], r[530], c[530]);
FA FA_497(p[33][28], p[34][27], p[35][26], r[531], c[531]);
FA FA_498(p[36][25], p[37][24], p[38][23], r[532], c[532]);
FA FA_499(p[39][22], p[40][21], p[41][20], r[533], c[533]);
FA FA_500(p[42][19], p[43][18], p[44][17], r[534], c[534]);
FA FA_501(p[26][36], p[27][35], p[28][34], r[535], c[535]);
FA FA_502(p[29][33], p[30][32], p[31][31], r[536], c[536]);
FA FA_503(p[32][30], p[33][29], p[34][28], r[537], c[537]);
FA FA_504(p[35][27], p[36][26], p[37][25], r[538], c[538]);
FA FA_505(p[38][24], p[39][23], p[40][22], r[539], c[539]);
FA FA_506(p[41][21], p[42][20], p[43][19], r[540], c[540]);
FA FA_507(p[44][18], p[45][17], p[46][16], r[541], c[541]);
FA FA_508(p[24][39], p[25][38], p[26][37], r[542], c[542]);
FA FA_509(p[27][36], p[28][35], p[29][34], r[543], c[543]);
FA FA_510(p[30][33], p[31][32], p[32][31], r[544], c[544]);
FA FA_511(p[33][30], p[34][29], p[35][28], r[545], c[545]);
FA FA_512(p[36][27], p[37][26], p[38][25], r[546], c[546]);
FA FA_513(p[39][24], p[40][23], p[41][22], r[547], c[547]);
FA FA_514(p[42][21], p[43][20], p[44][19], r[548], c[548]);
FA FA_515(c[3], r[4], c[297], r[549], c[549]);
FA FA_516(c[4], r[5], c[298], r[550], c[550]);
HA HA_34(r[299], c[549], r[551], c[551]);
FA FA_517(r[6], r[7], c[299], r[552], c[552]);
FA FA_518(p[6][1], p[7][0], c[6], r[553], c[553]);
HA HA_35(c[7], r[8], r[554], c[554]);
FA FA_519(p[6][2], p[7][1], p[8][0], r[555], c[555]);
FA FA_520(p[8][1], p[9][0], c[9], r[556], c[556]);
HA HA_36(r[10], r[11], r[557], c[557]);
FA FA_521(p[9][1], p[10][0], c[10], r[558], c[558]);
FA FA_522(p[11][0], c[12], c[13], r[559], c[559]);
FA FA_523(p[12][0], c[14], c[15], r[560], c[560]);
FA FA_524(c[17], c[18], r[19], r[561], c[561]);
FA FA_525(p[14][0], c[19], c[20], r[562], c[562]);
FA FA_526(r[21], r[22], r[23], r[563], c[563]);
FA FA_527(p[14][1], p[15][0], c[21], r[564], c[564]);
FA FA_528(c[22], c[23], r[24], r[565], c[565]);
HA HA_37(r[25], c[311], r[566], c[566]);
FA FA_529(p[12][4], p[13][3], p[14][2], r[567], c[567]);
FA FA_530(p[15][1], p[16][0], c[24], r[568], c[568]);
HA HA_38(c[25], r[26], r[569], c[569]);
FA FA_531(p[16][1], p[17][0], c[26], r[570], c[570]);
FA FA_532(c[27], r[28], r[29], r[571], c[571]);
FA FA_533(p[15][3], p[16][2], p[17][1], r[572], c[572]);
FA FA_534(p[18][0], c[28], c[29], r[573], c[573]);
HA HA_39(c[30], r[31], r[574], c[574]);
FA FA_535(p[17][2], p[18][1], p[19][0], r[575], c[575]);
FA FA_536(c[31], c[32], c[33], r[576], c[576]);
HA HA_40(r[34], r[35], r[577], c[577]);
FA FA_537(p[18][2], p[19][1], p[20][0], r[578], c[578]);
FA FA_538(c[34], c[35], c[36], r[579], c[579]);
FA FA_539(p[18][3], p[19][2], p[20][1], r[580], c[580]);
FA FA_540(p[21][0], c[38], c[39], r[581], c[581]);
FA FA_541(p[20][2], p[21][1], p[22][0], r[582], c[582]);
FA FA_542(c[41], c[42], c[43], r[583], c[583]);
FA FA_543(p[18][5], p[19][4], p[20][3], r[584], c[584]);
FA FA_544(p[21][2], p[22][1], p[23][0], r[585], c[585]);
FA FA_545(c[44], c[45], c[46], r[586], c[586]);
FA FA_546(p[18][6], p[19][5], p[20][4], r[587], c[587]);
FA FA_547(p[21][3], p[22][2], p[23][1], r[588], c[588]);
FA FA_548(p[24][0], c[48], c[49], r[589], c[589]);
FA FA_549(p[20][5], p[21][4], p[22][3], r[590], c[590]);
FA FA_550(p[23][2], p[24][1], p[25][0], r[591], c[591]);
FA FA_551(c[51], c[52], c[53], r[592], c[592]);
FA FA_552(p[23][3], p[24][2], p[25][1], r[593], c[593]);
FA FA_553(p[26][0], c[54], c[55], r[594], c[594]);
FA FA_554(c[56], c[57], r[58], r[595], c[595]);
FA FA_555(p[23][4], p[24][3], p[25][2], r[596], c[596]);
FA FA_556(p[26][1], p[27][0], c[58], r[597], c[597]);
FA FA_557(c[59], c[60], c[61], r[598], c[598]);
FA FA_558(p[23][5], p[24][4], p[25][3], r[599], c[599]);
FA FA_559(p[26][2], p[27][1], p[28][0], r[600], c[600]);
FA FA_560(c[62], c[63], c[64], r[601], c[601]);
FA FA_561(p[24][5], p[25][4], p[26][3], r[602], c[602]);
FA FA_562(p[27][2], p[28][1], p[29][0], r[603], c[603]);
FA FA_563(c[67], c[68], c[69], r[604], c[604]);
FA FA_564(p[26][4], p[27][3], p[28][2], r[605], c[605]);
FA FA_565(p[29][1], p[30][0], c[71], r[606], c[606]);
FA FA_566(c[72], c[73], c[74], r[607], c[607]);
FA FA_567(p[24][7], p[25][6], p[26][5], r[608], c[608]);
FA FA_568(p[27][4], p[28][3], p[29][2], r[609], c[609]);
FA FA_569(p[30][1], p[31][0], c[75], r[610], c[610]);
FA FA_570(p[24][8], p[25][7], p[26][6], r[611], c[611]);
FA FA_571(p[27][5], p[28][4], p[29][3], r[612], c[612]);
FA FA_572(p[30][2], p[31][1], p[32][0], r[613], c[613]);
FA FA_573(p[26][7], p[27][6], p[28][5], r[614], c[614]);
FA FA_574(p[29][4], p[30][3], p[31][2], r[615], c[615]);
FA FA_575(p[32][1], p[33][0], c[84], r[616], c[616]);
FA FA_576(p[27][7], p[28][6], p[29][5], r[617], c[617]);
FA FA_577(p[30][4], p[31][3], p[32][2], r[618], c[618]);
FA FA_578(p[33][1], p[34][0], c[88], r[619], c[619]);
HA HA_41(c[89], c[90], r[620], c[620]);
FA FA_579(p[29][6], p[30][5], p[31][4], r[621], c[621]);
FA FA_580(p[32][3], p[33][2], p[34][1], r[622], c[622]);
FA FA_581(p[35][0], c[93], c[94], r[623], c[623]);
FA FA_582(c[95], c[96], c[97], r[624], c[624]);
FA FA_583(p[27][9], p[28][8], p[29][7], r[625], c[625]);
FA FA_584(p[30][6], p[31][5], p[32][4], r[626], c[626]);
FA FA_585(p[33][3], p[34][2], p[35][1], r[627], c[627]);
FA FA_586(p[36][0], c[98], c[99], r[628], c[628]);
FA FA_587(p[27][10], p[28][9], p[29][8], r[629], c[629]);
FA FA_588(p[30][7], p[31][6], p[32][5], r[630], c[630]);
FA FA_589(p[33][4], p[34][3], p[35][2], r[631], c[631]);
FA FA_590(p[36][1], p[37][0], c[104], r[632], c[632]);
FA FA_591(p[29][9], p[30][8], p[31][7], r[633], c[633]);
FA FA_592(p[32][6], p[33][5], p[34][4], r[634], c[634]);
FA FA_593(p[35][3], p[36][2], p[37][1], r[635], c[635]);
FA FA_594(p[38][0], c[109], c[110], r[636], c[636]);
FA FA_595(p[30][9], p[31][8], p[32][7], r[637], c[637]);
FA FA_596(p[33][6], p[34][5], p[35][4], r[638], c[638]);
FA FA_597(p[36][3], p[37][2], p[38][1], r[639], c[639]);
FA FA_598(p[39][0], c[114], c[115], r[640], c[640]);
FA FA_599(p[32][8], p[33][7], p[34][6], r[641], c[641]);
FA FA_600(p[35][5], p[36][4], p[37][3], r[642], c[642]);
FA FA_601(p[38][2], p[39][1], p[40][0], r[643], c[643]);
FA FA_602(c[120], c[121], c[122], r[644], c[644]);
FA FA_603(p[32][9], p[33][8], p[34][7], r[645], c[645]);
FA FA_604(p[35][6], p[36][5], p[37][4], r[646], c[646]);
FA FA_605(p[38][3], p[39][2], p[40][1], r[647], c[647]);
FA FA_606(p[41][0], c[125], c[126], r[648], c[648]);
FA FA_607(p[33][9], p[34][8], p[35][7], r[649], c[649]);
FA FA_608(p[36][6], p[37][5], p[38][4], r[650], c[650]);
FA FA_609(p[39][3], p[40][2], p[41][1], r[651], c[651]);
FA FA_610(p[42][0], c[130], c[131], r[652], c[652]);
FA FA_611(p[35][8], p[36][7], p[37][6], r[653], c[653]);
FA FA_612(p[38][5], p[39][4], p[40][3], r[654], c[654]);
FA FA_613(p[41][2], p[42][1], p[43][0], r[655], c[655]);
FA FA_614(c[136], c[137], c[138], r[656], c[656]);
FA FA_615(p[33][11], p[34][10], p[35][9], r[657], c[657]);
FA FA_616(p[36][8], p[37][7], p[38][6], r[658], c[658]);
FA FA_617(p[39][5], p[40][4], p[41][3], r[659], c[659]);
FA FA_618(p[42][2], p[43][1], p[44][0], r[660], c[660]);
FA FA_619(c[142], c[143], c[144], r[661], c[661]);
FA FA_620(p[33][12], p[34][11], p[35][10], r[662], c[662]);
FA FA_621(p[36][9], p[37][8], p[38][7], r[663], c[663]);
FA FA_622(p[39][6], p[40][5], p[41][4], r[664], c[664]);
FA FA_623(p[42][3], p[43][2], p[44][1], r[665], c[665]);
FA FA_624(p[45][0], c[149], c[150], r[666], c[666]);
FA FA_625(p[35][11], p[36][10], p[37][9], r[667], c[667]);
FA FA_626(p[38][8], p[39][7], p[40][6], r[668], c[668]);
FA FA_627(p[41][5], p[42][4], p[43][3], r[669], c[669]);
FA FA_628(p[44][2], p[45][1], p[46][0], r[670], c[670]);
FA FA_629(c[155], c[156], c[157], r[671], c[671]);
FA FA_630(p[36][11], p[37][10], p[38][9], r[672], c[672]);
FA FA_631(p[39][8], p[40][7], p[41][6], r[673], c[673]);
FA FA_632(p[42][5], p[43][4], p[44][3], r[674], c[674]);
FA FA_633(p[45][2], p[46][1], p[47][0], r[675], c[675]);
FA FA_634(c[161], c[162], c[163], r[676], c[676]);
HA HA_42(c[164], c[165], r[677], c[677]);
FA FA_635(p[36][12], p[37][11], p[38][10], r[678], c[678]);
FA FA_636(p[39][9], p[40][8], p[41][7], r[679], c[679]);
FA FA_637(p[42][6], p[43][5], p[44][4], r[680], c[680]);
FA FA_638(p[45][3], p[46][2], p[47][1], r[681], c[681]);
FA FA_639(p[48][0], c[168], c[169], r[682], c[682]);
FA FA_640(p[38][11], p[39][10], p[40][9], r[683], c[683]);
FA FA_641(p[41][8], p[42][7], p[43][6], r[684], c[684]);
FA FA_642(p[44][5], p[45][4], p[46][3], r[685], c[685]);
FA FA_643(p[47][2], p[48][1], p[49][0], r[686], c[686]);
FA FA_644(c[174], c[175], c[176], r[687], c[687]);
FA FA_645(p[41][9], p[42][8], p[43][7], r[688], c[688]);
FA FA_646(p[44][6], p[45][5], p[46][4], r[689], c[689]);
FA FA_647(p[47][3], p[48][2], p[49][1], r[690], c[690]);
FA FA_648(p[50][0], c[180], c[181], r[691], c[691]);
FA FA_649(c[182], c[183], c[184], r[692], c[692]);
FA FA_650(p[41][10], p[42][9], p[43][8], r[693], c[693]);
FA FA_651(p[44][7], p[45][6], p[46][5], r[694], c[694]);
FA FA_652(p[47][4], p[48][3], p[49][2], r[695], c[695]);
FA FA_653(p[50][1], p[51][0], c[187], r[696], c[696]);
FA FA_654(c[188], c[189], c[190], r[697], c[697]);
HA HA_43(c[191], c[192], r[698], c[698]);
FA FA_655(p[41][11], p[42][10], p[43][9], r[699], c[699]);
FA FA_656(p[44][8], p[45][7], p[46][6], r[700], c[700]);
FA FA_657(p[47][5], p[48][4], p[49][3], r[701], c[701]);
FA FA_658(p[50][2], p[51][1], p[52][0], r[702], c[702]);
FA FA_659(c[194], c[195], c[196], r[703], c[703]);
FA FA_660(p[39][14], p[40][13], p[41][12], r[704], c[704]);
FA FA_661(p[42][11], p[43][10], p[44][9], r[705], c[705]);
FA FA_662(p[45][8], p[46][7], p[47][6], r[706], c[706]);
FA FA_663(p[48][5], p[49][4], p[50][3], r[707], c[707]);
FA FA_664(p[51][2], p[52][1], p[53][0], r[708], c[708]);
HA HA_44(c[202], c[203], r[709], c[709]);
FA FA_665(p[43][11], p[44][10], p[45][9], r[710], c[710]);
FA FA_666(p[46][8], p[47][7], p[48][6], r[711], c[711]);
FA FA_667(p[49][5], p[50][4], p[51][3], r[712], c[712]);
FA FA_668(p[52][2], p[53][1], p[54][0], r[713], c[713]);
FA FA_669(c[209], c[210], c[211], r[714], c[714]);
FA FA_670(p[42][13], p[43][12], p[44][11], r[715], c[715]);
FA FA_671(p[45][10], p[46][9], p[47][8], r[716], c[716]);
FA FA_672(p[48][7], p[49][6], p[50][5], r[717], c[717]);
FA FA_673(p[51][4], p[52][3], p[53][2], r[718], c[718]);
FA FA_674(p[54][1], p[55][0], c[216], r[719], c[719]);
FA FA_675(c[217], c[218], c[219], r[720], c[720]);
FA FA_676(p[42][14], p[43][13], p[44][12], r[721], c[721]);
FA FA_677(p[45][11], p[46][10], p[47][9], r[722], c[722]);
FA FA_678(p[48][8], p[49][7], p[50][6], r[723], c[723]);
FA FA_679(p[51][5], p[52][4], p[53][3], r[724], c[724]);
FA FA_680(p[54][2], p[55][1], p[56][0], r[725], c[725]);
FA FA_681(c[224], c[225], c[226], r[726], c[726]);
FA FA_682(p[44][13], p[45][12], p[46][11], r[727], c[727]);
FA FA_683(p[47][10], p[48][9], p[49][8], r[728], c[728]);
FA FA_684(p[50][7], p[51][6], p[52][5], r[729], c[729]);
FA FA_685(p[53][4], p[54][3], p[55][2], r[730], c[730]);
FA FA_686(p[56][1], p[57][0], c[231], r[731], c[731]);
FA FA_687(c[232], c[233], c[234], r[732], c[732]);
FA FA_688(p[45][13], p[46][12], p[47][11], r[733], c[733]);
FA FA_689(p[48][10], p[49][9], p[50][8], r[734], c[734]);
FA FA_690(p[51][7], p[52][6], p[53][5], r[735], c[735]);
FA FA_691(p[54][4], p[55][3], p[56][2], r[736], c[736]);
FA FA_692(p[57][1], p[58][0], c[238], r[737], c[737]);
FA FA_693(c[239], c[240], c[241], r[738], c[738]);
HA HA_45(c[242], c[243], r[739], c[739]);
FA FA_694(p[47][12], p[48][11], p[49][10], r[740], c[740]);
FA FA_695(p[50][9], p[51][8], p[52][7], r[741], c[741]);
FA FA_696(p[53][6], p[54][5], p[55][4], r[742], c[742]);
FA FA_697(p[56][3], p[57][2], p[58][1], r[743], c[743]);
FA FA_698(p[59][0], c[246], c[247], r[744], c[744]);
FA FA_699(c[248], c[249], c[250], r[745], c[745]);
FA FA_700(p[45][15], p[46][14], p[47][13], r[746], c[746]);
FA FA_701(p[48][12], p[49][11], p[50][10], r[747], c[747]);
FA FA_702(p[51][9], p[52][8], p[53][7], r[748], c[748]);
FA FA_703(p[54][6], p[55][5], p[56][4], r[749], c[749]);
FA FA_704(p[57][3], p[58][2], p[59][1], r[750], c[750]);
FA FA_705(p[60][0], c[254], c[255], r[751], c[751]);
HA HA_46(c[256], c[257], r[752], c[752]);
FA FA_706(p[45][16], p[46][15], p[47][14], r[753], c[753]);
FA FA_707(p[48][13], p[49][12], p[50][11], r[754], c[754]);
FA FA_708(p[51][10], p[52][9], p[53][8], r[755], c[755]);
FA FA_709(p[54][7], p[55][6], p[56][5], r[756], c[756]);
FA FA_710(p[57][4], p[58][3], p[59][2], r[757], c[757]);
FA FA_711(p[60][1], p[61][0], c[263], r[758], c[758]);
FA FA_712(p[47][15], p[48][14], p[49][13], r[759], c[759]);
FA FA_713(p[50][12], p[51][11], p[52][10], r[760], c[760]);
FA FA_714(p[53][9], p[54][8], p[55][7], r[761], c[761]);
FA FA_715(p[56][6], p[57][5], p[58][4], r[762], c[762]);
FA FA_716(p[59][3], p[60][2], p[61][1], r[763], c[763]);
FA FA_717(p[62][0], c[271], c[272], r[764], c[764]);
HA HA_47(c[273], c[274], r[765], c[765]);
FA FA_718(p[45][18], p[46][17], p[47][16], r[766], c[766]);
FA FA_719(p[48][15], p[49][14], p[50][13], r[767], c[767]);
FA FA_720(p[51][12], p[52][11], p[53][10], r[768], c[768]);
FA FA_721(p[54][9], p[55][8], p[56][7], r[769], c[769]);
FA FA_722(p[57][6], p[58][5], p[59][4], r[770], c[770]);
FA FA_723(p[60][3], p[61][2], p[62][1], r[771], c[771]);
FA FA_724(p[63][0], c[279], c[280], r[772], c[772]);
HA HA_48(r[298], r[549], r[773], c[773]);
FA FA_725(r[550], r[551], c[773], r[774], c[774]);
FA FA_726(r[300], c[550], c[551], r[775], c[775]);
HA HA_49(r[552], c[774], r[776], c[776]);
FA FA_727(c[300], r[301], c[552], r[777], c[777]);
FA FA_728(c[8], r[9], c[301], r[778], c[778]);
HA HA_50(r[302], c[553], r[779], c[779]);
FA FA_729(c[302], r[303], c[555], r[780], c[780]);
FA FA_730(c[11], r[12], r[13], r[781], c[781]);
FA FA_731(r[14], r[15], r[16], r[782], c[782]);
HA HA_51(c[304], r[305], r[783], c[783]);
FA FA_732(c[16], r[17], r[18], r[784], c[784]);
FA FA_733(r[20], c[306], c[307], r[785], c[785]);
FA FA_734(c[308], c[309], c[310], r[786], c[786]);
FA FA_735(c[312], r[313], r[314], r[787], c[787]);
FA FA_736(r[27], c[313], c[314], r[788], c[788]);
FA FA_737(c[315], r[316], r[317], r[789], c[789]);
FA FA_738(r[30], c[316], c[317], r[790], c[790]);
FA FA_739(r[318], r[319], r[320], r[791], c[791]);
FA FA_740(r[32], r[33], c[318], r[792], c[792]);
FA FA_741(c[319], c[320], r[321], r[793], c[793]);
HA HA_52(r[322], c[570], r[794], c[794]);
FA FA_742(r[36], r[37], c[321], r[795], c[795]);
FA FA_743(c[322], r[323], r[324], r[796], c[796]);
FA FA_744(c[37], r[38], r[39], r[797], c[797]);
FA FA_745(r[40], c[323], c[324], r[798], c[798]);
FA FA_746(c[40], r[41], r[42], r[799], c[799]);
FA FA_747(r[43], c[325], c[326], r[800], c[800]);
FA FA_748(r[44], r[45], r[46], r[801], c[801]);
FA FA_749(r[47], c[328], c[329], r[802], c[802]);
FA FA_750(c[47], r[48], r[49], r[803], c[803]);
FA FA_751(r[50], c[331], c[332], r[804], c[804]);
HA HA_53(c[333], r[334], r[805], c[805]);
FA FA_752(c[50], r[51], r[52], r[806], c[806]);
FA FA_753(r[53], c[334], c[335], r[807], c[807]);
FA FA_754(r[54], r[55], r[56], r[808], c[808]);
FA FA_755(r[57], c[337], c[338], r[809], c[809]);
FA FA_756(r[59], r[60], r[61], r[810], c[810]);
FA FA_757(c[340], c[341], c[342], r[811], c[811]);
FA FA_758(r[62], r[63], r[64], r[812], c[812]);
FA FA_759(r[65], r[66], c[343], r[813], c[813]);
HA HA_54(c[344], c[345], r[814], c[814]);
FA FA_760(c[65], c[66], r[67], r[815], c[815]);
FA FA_761(r[68], r[69], r[70], r[816], c[816]);
FA FA_762(c[347], c[348], c[349], r[817], c[817]);
FA FA_763(c[70], r[71], r[72], r[818], c[818]);
FA FA_764(r[73], r[74], c[350], r[819], c[819]);
FA FA_765(c[351], c[352], c[353], r[820], c[820]);
FA FA_766(r[75], r[76], r[77], r[821], c[821]);
FA FA_767(r[78], r[79], c[354], r[822], c[822]);
FA FA_768(c[355], c[356], c[357], r[823], c[823]);
FA FA_769(c[76], c[77], c[78], r[824], c[824]);
FA FA_770(c[79], r[80], r[81], r[825], c[825]);
FA FA_771(r[82], r[83], c[358], r[826], c[826]);
FA FA_772(c[80], c[81], c[82], r[827], c[827]);
FA FA_773(c[83], r[84], r[85], r[828], c[828]);
FA FA_774(r[86], r[87], c[362], r[829], c[829]);
FA FA_775(c[85], c[86], c[87], r[830], c[830]);
FA FA_776(r[88], r[89], r[90], r[831], c[831]);
FA FA_777(r[91], r[92], c[366], r[832], c[832]);
FA FA_778(c[91], c[92], r[93], r[833], c[833]);
FA FA_779(r[94], r[95], r[96], r[834], c[834]);
FA FA_780(r[97], c[370], c[371], r[835], c[835]);
FA FA_781(r[98], r[99], r[100], r[836], c[836]);
FA FA_782(r[101], r[102], r[103], r[837], c[837]);
FA FA_783(c[374], c[375], c[376], r[838], c[838]);
FA FA_784(c[100], c[101], c[102], r[839], c[839]);
FA FA_785(c[103], r[104], r[105], r[840], c[840]);
FA FA_786(r[106], r[107], r[108], r[841], c[841]);
FA FA_787(c[105], c[106], c[107], r[842], c[842]);
FA FA_788(c[108], r[109], r[110], r[843], c[843]);
FA FA_789(r[111], r[112], r[113], r[844], c[844]);
FA FA_790(c[111], c[112], c[113], r[845], c[845]);
FA FA_791(r[114], r[115], r[116], r[846], c[846]);
FA FA_792(r[117], r[118], r[119], r[847], c[847]);
FA FA_793(c[116], c[117], c[118], r[848], c[848]);
FA FA_794(c[119], r[120], r[121], r[849], c[849]);
FA FA_795(r[122], r[123], r[124], r[850], c[850]);
HA HA_55(c[390], c[391], r[851], c[851]);
FA FA_796(c[123], c[124], r[125], r[852], c[852]);
FA FA_797(r[126], r[127], r[128], r[853], c[853]);
FA FA_798(r[129], c[394], c[395], r[854], c[854]);
FA FA_799(c[396], c[397], c[398], r[855], c[855]);
FA FA_800(c[127], c[128], c[129], r[856], c[856]);
FA FA_801(r[130], r[131], r[132], r[857], c[857]);
FA FA_802(r[133], r[134], r[135], r[858], c[858]);
FA FA_803(c[399], c[400], c[401], r[859], c[859]);
HA HA_56(c[402], c[403], r[860], c[860]);
FA FA_804(c[132], c[133], c[134], r[861], c[861]);
FA FA_805(c[135], r[136], r[137], r[862], c[862]);
FA FA_806(r[138], r[139], r[140], r[863], c[863]);
FA FA_807(r[141], c[405], c[406], r[864], c[864]);
FA FA_808(c[139], c[140], c[141], r[865], c[865]);
FA FA_809(r[142], r[143], r[144], r[866], c[866]);
FA FA_810(r[145], r[146], r[147], r[867], c[867]);
FA FA_811(r[148], c[410], c[411], r[868], c[868]);
HA HA_57(c[412], c[413], r[869], c[869]);
FA FA_812(c[145], c[146], c[147], r[870], c[870]);
FA FA_813(c[148], r[149], r[150], r[871], c[871]);
FA FA_814(r[151], r[152], r[153], r[872], c[872]);
FA FA_815(r[154], c[415], c[416], r[873], c[873]);
FA FA_816(c[151], c[152], c[153], r[874], c[874]);
FA FA_817(c[154], r[155], r[156], r[875], c[875]);
FA FA_818(r[157], r[158], r[159], r[876], c[876]);
FA FA_819(r[160], c[420], c[421], r[877], c[877]);
FA FA_820(c[158], c[159], c[160], r[878], c[878]);
FA FA_821(r[161], r[162], r[163], r[879], c[879]);
FA FA_822(r[164], r[165], r[166], r[880], c[880]);
FA FA_823(r[167], c[425], c[426], r[881], c[881]);
FA FA_824(c[166], c[167], r[168], r[882], c[882]);
FA FA_825(r[169], r[170], r[171], r[883], c[883]);
FA FA_826(r[172], r[173], c[430], r[884], c[884]);
FA FA_827(c[431], c[432], c[433], r[885], c[885]);
FA FA_828(c[170], c[171], c[172], r[886], c[886]);
FA FA_829(c[173], r[174], r[175], r[887], c[887]);
FA FA_830(r[176], r[177], r[178], r[888], c[888]);
FA FA_831(r[179], c[435], c[436], r[889], c[889]);
FA FA_832(c[177], c[178], c[179], r[890], c[890]);
FA FA_833(r[180], r[181], r[182], r[891], c[891]);
FA FA_834(r[183], r[184], r[185], r[892], c[892]);
FA FA_835(r[186], c[441], c[442], r[893], c[893]);
FA FA_836(c[185], c[186], r[187], r[894], c[894]);
FA FA_837(r[188], r[189], r[190], r[895], c[895]);
FA FA_838(r[191], r[192], r[193], r[896], c[896]);
FA FA_839(c[447], c[448], c[449], r[897], c[897]);
FA FA_840(c[193], r[194], r[195], r[898], c[898]);
FA FA_841(r[196], r[197], r[198], r[899], c[899]);
FA FA_842(r[199], r[200], r[201], r[900], c[900]);
FA FA_843(c[453], c[454], c[455], r[901], c[901]);
FA FA_844(c[197], c[198], c[199], r[902], c[902]);
FA FA_845(c[200], c[201], r[202], r[903], c[903]);
FA FA_846(r[203], r[204], r[205], r[904], c[904]);
FA FA_847(r[206], r[207], r[208], r[905], c[905]);
FA FA_848(c[460], c[461], c[462], r[906], c[906]);
FA FA_849(c[204], c[205], c[206], r[907], c[907]);
FA FA_850(c[207], c[208], r[209], r[908], c[908]);
FA FA_851(r[210], r[211], r[212], r[909], c[909]);
FA FA_852(r[213], r[214], r[215], r[910], c[910]);
FA FA_853(c[466], c[467], c[468], r[911], c[911]);
HA HA_58(c[469], c[470], r[912], c[912]);
FA FA_854(c[212], c[213], c[214], r[913], c[913]);
FA FA_855(c[215], r[216], r[217], r[914], c[914]);
FA FA_856(r[218], r[219], r[220], r[915], c[915]);
FA FA_857(r[221], r[222], r[223], r[916], c[916]);
FA FA_858(c[473], c[474], c[475], r[917], c[917]);
FA FA_859(c[220], c[221], c[222], r[918], c[918]);
FA FA_860(c[223], r[224], r[225], r[919], c[919]);
FA FA_861(r[226], r[227], r[228], r[920], c[920]);
FA FA_862(r[229], r[230], c[479], r[921], c[921]);
FA FA_863(c[480], c[481], c[482], r[922], c[922]);
HA HA_59(c[483], c[484], r[923], c[923]);
FA FA_864(c[227], c[228], c[229], r[924], c[924]);
FA FA_865(c[230], r[231], r[232], r[925], c[925]);
FA FA_866(r[233], r[234], r[235], r[926], c[926]);
FA FA_867(r[236], r[237], c[486], r[927], c[927]);
FA FA_868(c[487], c[488], c[489], r[928], c[928]);
FA FA_869(c[235], c[236], c[237], r[929], c[929]);
FA FA_870(r[238], r[239], r[240], r[930], c[930]);
FA FA_871(r[241], r[242], r[243], r[931], c[931]);
FA FA_872(r[244], r[245], c[493], r[932], c[932]);
FA FA_873(c[494], c[495], c[496], r[933], c[933]);
FA FA_874(c[244], c[245], r[246], r[934], c[934]);
FA FA_875(r[247], r[248], r[249], r[935], c[935]);
FA FA_876(r[250], r[251], r[252], r[936], c[936]);
FA FA_877(r[253], c[500], c[501], r[937], c[937]);
FA FA_878(c[502], c[503], c[504], r[938], c[938]);
FA FA_879(c[251], c[252], c[253], r[939], c[939]);
FA FA_880(r[254], r[255], r[256], r[940], c[940]);
FA FA_881(r[257], r[258], r[259], r[941], c[941]);
FA FA_882(r[260], r[261], r[262], r[942], c[942]);
FA FA_883(c[507], c[508], c[509], r[943], c[943]);
HA HA_60(c[510], c[511], r[944], c[944]);
FA FA_884(c[258], c[259], c[260], r[945], c[945]);
FA FA_885(c[261], c[262], r[263], r[946], c[946]);
FA FA_886(r[264], r[265], r[266], r[947], c[947]);
FA FA_887(r[267], r[268], r[269], r[948], c[948]);
FA FA_888(r[270], c[514], c[515], r[949], c[949]);
FA FA_889(c[264], c[265], c[266], r[950], c[950]);
FA FA_890(c[267], c[268], c[269], r[951], c[951]);
FA FA_891(c[270], r[271], r[272], r[952], c[952]);
FA FA_892(r[273], r[274], r[275], r[953], c[953]);
FA FA_893(r[276], r[277], r[278], r[954], c[954]);
HA HA_61(c[521], c[522], r[955], c[955]);
FA FA_894(c[275], c[276], c[277], r[956], c[956]);
FA FA_895(c[278], r[279], r[280], r[957], c[957]);
FA FA_896(r[281], r[282], r[283], r[958], c[958]);
FA FA_897(r[284], r[285], r[286], r[959], c[959]);
FA FA_898(r[287], c[528], c[529], r[960], c[960]);
FA FA_899(c[281], c[282], c[283], r[961], c[961]);
FA FA_900(c[284], c[285], c[286], r[962], c[962]);
FA FA_901(c[287], r[288], r[289], r[963], c[963]);
FA FA_902(r[290], r[291], r[292], r[964], c[964]);
FA FA_903(r[293], r[294], r[295], r[965], c[965]);
FA FA_904(c[535], c[536], c[537], r[966], c[966]);
HA HA_62(r[775], r[776], r[967], c[967]);
FA FA_905(r[553], r[554], c[775], r[968], c[968]);
FA FA_906(c[554], r[555], c[777], r[969], c[969]);
FA FA_907(r[556], r[557], c[778], r[970], c[970]);
FA FA_908(c[303], r[304], c[556], r[971], c[971]);
HA HA_63(c[557], r[558], r[972], c[972]);
FA FA_909(c[558], r[559], c[781], r[973], c[973]);
FA FA_910(c[305], r[306], r[307], r[974], c[974]);
FA FA_911(r[308], r[309], r[310], r[975], c[975]);
HA HA_64(c[560], r[561], r[976], c[976]);
FA FA_912(r[311], r[312], c[561], r[977], c[977]);
FA FA_913(r[315], c[562], c[563], r[978], c[978]);
FA FA_914(c[564], c[565], c[566], r[979], c[979]);
FA FA_915(c[567], c[568], c[569], r[980], c[980]);
FA FA_916(c[571], r[572], r[573], r[981], c[981]);
FA FA_917(c[572], c[573], c[574], r[982], c[982]);
FA FA_918(r[575], r[576], r[577], r[983], c[983]);
FA FA_919(r[325], r[326], r[327], r[984], c[984]);
FA FA_920(c[575], c[576], c[577], r[985], c[985]);
HA HA_65(r[578], r[579], r[986], c[986]);
FA FA_921(c[327], r[328], r[329], r[987], c[987]);
FA FA_922(r[330], c[578], c[579], r[988], c[988]);
FA FA_923(c[330], r[331], r[332], r[989], c[989]);
FA FA_924(r[333], c[580], c[581], r[990], c[990]);
HA HA_66(r[582], r[583], r[991], c[991]);
FA FA_925(r[335], r[336], c[582], r[992], c[992]);
FA FA_926(c[583], r[584], r[585], r[993], c[993]);
FA FA_927(c[336], r[337], r[338], r[994], c[994]);
FA FA_928(r[339], c[584], c[585], r[995], c[995]);
HA HA_67(c[586], r[587], r[996], c[996]);
FA FA_929(c[339], r[340], r[341], r[997], c[997]);
FA FA_930(r[342], c[587], c[588], r[998], c[998]);
HA HA_68(c[589], r[590], r[999], c[999]);
FA FA_931(r[343], r[344], r[345], r[1000], c[1000]);
FA FA_932(r[346], c[590], c[591], r[1001], c[1001]);
HA HA_69(c[592], r[593], r[1002], c[1002]);
FA FA_933(c[346], r[347], r[348], r[1003], c[1003]);
FA FA_934(r[349], c[593], c[594], r[1004], c[1004]);
FA FA_935(r[350], r[351], r[352], r[1005], c[1005]);
FA FA_936(r[353], c[596], c[597], r[1006], c[1006]);
FA FA_937(r[354], r[355], r[356], r[1007], c[1007]);
FA FA_938(r[357], c[599], c[600], r[1008], c[1008]);
FA FA_939(r[358], r[359], r[360], r[1009], c[1009]);
FA FA_940(r[361], c[602], c[603], r[1010], c[1010]);
FA FA_941(c[359], c[360], c[361], r[1011], c[1011]);
FA FA_942(r[362], r[363], r[364], r[1012], c[1012]);
FA FA_943(r[365], c[605], c[606], r[1013], c[1013]);
FA FA_944(c[363], c[364], c[365], r[1014], c[1014]);
FA FA_945(r[366], r[367], r[368], r[1015], c[1015]);
FA FA_946(r[369], c[608], c[609], r[1016], c[1016]);
FA FA_947(c[367], c[368], c[369], r[1017], c[1017]);
FA FA_948(r[370], r[371], r[372], r[1018], c[1018]);
FA FA_949(r[373], c[611], c[612], r[1019], c[1019]);
FA FA_950(c[372], c[373], r[374], r[1020], c[1020]);
FA FA_951(r[375], r[376], r[377], r[1021], c[1021]);
FA FA_952(c[614], c[615], c[616], r[1022], c[1022]);
FA FA_953(c[377], r[378], r[379], r[1023], c[1023]);
FA FA_954(r[380], r[381], c[617], r[1024], c[1024]);
FA FA_955(c[618], c[619], c[620], r[1025], c[1025]);
FA FA_956(c[378], c[379], c[380], r[1026], c[1026]);
FA FA_957(c[381], r[382], r[383], r[1027], c[1027]);
FA FA_958(r[384], r[385], c[621], r[1028], c[1028]);
FA FA_959(c[382], c[383], c[384], r[1029], c[1029]);
FA FA_960(c[385], r[386], r[387], r[1030], c[1030]);
FA FA_961(r[388], r[389], c[625], r[1031], c[1031]);
FA FA_962(c[386], c[387], c[388], r[1032], c[1032]);
FA FA_963(c[389], r[390], r[391], r[1033], c[1033]);
FA FA_964(r[392], r[393], c[629], r[1034], c[1034]);
FA FA_965(c[392], c[393], r[394], r[1035], c[1035]);
FA FA_966(r[395], r[396], r[397], r[1036], c[1036]);
FA FA_967(r[398], c[633], c[634], r[1037], c[1037]);
FA FA_968(r[399], r[400], r[401], r[1038], c[1038]);
FA FA_969(r[402], r[403], r[404], r[1039], c[1039]);
FA FA_970(c[637], c[638], c[639], r[1040], c[1040]);
FA FA_971(c[404], r[405], r[406], r[1041], c[1041]);
FA FA_972(r[407], r[408], r[409], r[1042], c[1042]);
FA FA_973(c[641], c[642], c[643], r[1043], c[1043]);
HA HA_70(c[644], r[645], r[1044], c[1044]);
FA FA_974(c[407], c[408], c[409], r[1045], c[1045]);
FA FA_975(r[410], r[411], r[412], r[1046], c[1046]);
FA FA_976(r[413], r[414], c[645], r[1047], c[1047]);
HA HA_71(c[646], c[647], r[1048], c[1048]);
FA FA_977(c[414], r[415], r[416], r[1049], c[1049]);
FA FA_978(r[417], r[418], r[419], r[1050], c[1050]);
FA FA_979(c[649], c[650], c[651], r[1051], c[1051]);
FA FA_980(c[417], c[418], c[419], r[1052], c[1052]);
FA FA_981(r[420], r[421], r[422], r[1053], c[1053]);
FA FA_982(r[423], r[424], c[653], r[1054], c[1054]);
HA HA_72(c[654], c[655], r[1055], c[1055]);
FA FA_983(c[422], c[423], c[424], r[1056], c[1056]);
FA FA_984(r[425], r[426], r[427], r[1057], c[1057]);
FA FA_985(r[428], r[429], c[657], r[1058], c[1058]);
FA FA_986(c[658], c[659], c[660], r[1059], c[1059]);
FA FA_987(c[427], c[428], c[429], r[1060], c[1060]);
FA FA_988(r[430], r[431], r[432], r[1061], c[1061]);
FA FA_989(r[433], r[434], c[662], r[1062], c[1062]);
FA FA_990(c[663], c[664], c[665], r[1063], c[1063]);
FA FA_991(c[434], r[435], r[436], r[1064], c[1064]);
FA FA_992(r[437], r[438], r[439], r[1065], c[1065]);
FA FA_993(r[440], c[667], c[668], r[1066], c[1066]);
FA FA_994(c[669], c[670], c[671], r[1067], c[1067]);
FA FA_995(c[437], c[438], c[439], r[1068], c[1068]);
FA FA_996(c[440], r[441], r[442], r[1069], c[1069]);
FA FA_997(r[443], r[444], r[445], r[1070], c[1070]);
FA FA_998(r[446], c[672], c[673], r[1071], c[1071]);
FA FA_999(c[443], c[444], c[445], r[1072], c[1072]);
FA FA_1000(c[446], r[447], r[448], r[1073], c[1073]);
FA FA_1001(r[449], r[450], r[451], r[1074], c[1074]);
FA FA_1002(r[452], c[678], c[679], r[1075], c[1075]);
HA HA_73(c[680], c[681], r[1076], c[1076]);
FA FA_1003(c[450], c[451], c[452], r[1077], c[1077]);
FA FA_1004(r[453], r[454], r[455], r[1078], c[1078]);
FA FA_1005(r[456], r[457], r[458], r[1079], c[1079]);
FA FA_1006(r[459], c[683], c[684], r[1080], c[1080]);
FA FA_1007(c[456], c[457], c[458], r[1081], c[1081]);
FA FA_1008(c[459], r[460], r[461], r[1082], c[1082]);
FA FA_1009(r[462], r[463], r[464], r[1083], c[1083]);
FA FA_1010(r[465], c[688], c[689], r[1084], c[1084]);
FA FA_1011(c[463], c[464], c[465], r[1085], c[1085]);
FA FA_1012(r[466], r[467], r[468], r[1086], c[1086]);
FA FA_1013(r[469], r[470], r[471], r[1087], c[1087]);
FA FA_1014(r[472], c[693], c[694], r[1088], c[1088]);
FA FA_1015(c[471], c[472], r[473], r[1089], c[1089]);
FA FA_1016(r[474], r[475], r[476], r[1090], c[1090]);
FA FA_1017(r[477], r[478], c[699], r[1091], c[1091]);
FA FA_1018(c[700], c[701], c[702], r[1092], c[1092]);
FA FA_1019(c[476], c[477], c[478], r[1093], c[1093]);
FA FA_1020(r[479], r[480], r[481], r[1094], c[1094]);
FA FA_1021(r[482], r[483], r[484], r[1095], c[1095]);
FA FA_1022(r[485], c[704], c[705], r[1096], c[1096]);
FA FA_1023(c[485], r[486], r[487], r[1097], c[1097]);
FA FA_1024(r[488], r[489], r[490], r[1098], c[1098]);
FA FA_1025(r[491], r[492], c[710], r[1099], c[1099]);
FA FA_1026(c[711], c[712], c[713], r[1100], c[1100]);
FA FA_1027(c[490], c[491], c[492], r[1101], c[1101]);
FA FA_1028(r[493], r[494], r[495], r[1102], c[1102]);
FA FA_1029(r[496], r[497], r[498], r[1103], c[1103]);
FA FA_1030(r[499], c[715], c[716], r[1104], c[1104]);
FA FA_1031(c[497], c[498], c[499], r[1105], c[1105]);
FA FA_1032(r[500], r[501], r[502], r[1106], c[1106]);
FA FA_1033(r[503], r[504], r[505], r[1107], c[1107]);
FA FA_1034(r[506], c[721], c[722], r[1108], c[1108]);
FA FA_1035(c[505], c[506], r[507], r[1109], c[1109]);
FA FA_1036(r[508], r[509], r[510], r[1110], c[1110]);
FA FA_1037(r[511], r[512], r[513], r[1111], c[1111]);
FA FA_1038(c[727], c[728], c[729], r[1112], c[1112]);
FA FA_1039(c[512], c[513], r[514], r[1113], c[1113]);
FA FA_1040(r[515], r[516], r[517], r[1114], c[1114]);
FA FA_1041(r[518], r[519], r[520], r[1115], c[1115]);
FA FA_1042(c[733], c[734], c[735], r[1116], c[1116]);
FA FA_1043(c[516], c[517], c[518], r[1117], c[1117]);
FA FA_1044(c[519], c[520], r[521], r[1118], c[1118]);
FA FA_1045(r[522], r[523], r[524], r[1119], c[1119]);
FA FA_1046(r[525], r[526], r[527], r[1120], c[1120]);
FA FA_1047(c[740], c[741], c[742], r[1121], c[1121]);
FA FA_1048(c[523], c[524], c[525], r[1122], c[1122]);
FA FA_1049(c[526], c[527], r[528], r[1123], c[1123]);
FA FA_1050(r[529], r[530], r[531], r[1124], c[1124]);
FA FA_1051(r[532], r[533], r[534], r[1125], c[1125]);
FA FA_1052(c[746], c[747], c[748], r[1126], c[1126]);
HA HA_74(c[749], c[750], r[1127], c[1127]);
FA FA_1053(c[530], c[531], c[532], r[1128], c[1128]);
FA FA_1054(c[533], c[534], r[535], r[1129], c[1129]);
FA FA_1055(r[536], r[537], r[538], r[1130], c[1130]);
FA FA_1056(r[539], r[540], r[541], r[1131], c[1131]);
FA FA_1057(c[753], c[754], c[755], r[1132], c[1132]);
FA FA_1058(c[538], c[539], c[540], r[1133], c[1133]);
FA FA_1059(c[541], r[542], r[543], r[1134], c[1134]);
FA FA_1060(r[544], r[545], r[546], r[1135], c[1135]);
FA FA_1061(r[547], r[548], c[759], r[1136], c[1136]);
FA FA_1062(c[760], c[761], c[762], r[1137], c[1137]);
HA HA_75(c[763], c[764], r[1138], c[1138]);
FA FA_1063(c[776], r[777], c[967], r[1139], c[1139]);
FA FA_1064(r[778], r[779], c[968], r[1140], c[1140]);
HA HA_76(r[969], c[1139], r[1141], c[1141]);
FA FA_1065(c[779], r[780], c[969], r[1142], c[1142]);
FA FA_1066(c[780], r[781], c[970], r[1143], c[1143]);
FA FA_1067(r[782], r[783], c[971], r[1144], c[1144]);
FA FA_1068(c[559], r[560], c[782], r[1145], c[1145]);
HA HA_77(c[783], r[784], r[1146], c[1146]);
FA FA_1069(c[784], r[785], c[974], r[1147], c[1147]);
FA FA_1070(r[562], r[563], c[785], r[1148], c[1148]);
HA HA_78(r[786], c[975], r[1149], c[1149]);
FA FA_1071(r[564], r[565], r[566], r[1150], c[1150]);
FA FA_1072(r[567], r[568], r[569], r[1151], c[1151]);
FA FA_1073(r[570], r[571], c[788], r[1152], c[1152]);
FA FA_1074(r[574], c[790], c[791], r[1153], c[1153]);
FA FA_1075(c[792], c[793], c[794], r[1154], c[1154]);
FA FA_1076(c[795], c[796], r[797], r[1155], c[1155]);
FA FA_1077(r[580], r[581], c[797], r[1156], c[1156]);
FA FA_1078(c[798], r[799], r[800], r[1157], c[1157]);
FA FA_1079(c[799], c[800], r[801], r[1158], c[1158]);
HA HA_79(r[802], c[987], r[1159], c[1159]);
FA FA_1080(r[586], c[801], c[802], r[1160], c[1160]);
FA FA_1081(r[803], r[804], r[805], r[1161], c[1161]);
FA FA_1082(r[588], r[589], c[803], r[1162], c[1162]);
FA FA_1083(c[804], c[805], r[806], r[1163], c[1163]);
HA HA_80(r[807], c[992], r[1164], c[1164]);
FA FA_1084(r[591], r[592], c[806], r[1165], c[1165]);
FA FA_1085(c[807], r[808], r[809], r[1166], c[1166]);
FA FA_1086(r[594], r[595], c[808], r[1167], c[1167]);
FA FA_1087(c[809], r[810], r[811], r[1168], c[1168]);
HA HA_81(c[997], c[998], r[1169], c[1169]);
FA FA_1088(c[595], r[596], r[597], r[1170], c[1170]);
FA FA_1089(r[598], c[810], c[811], r[1171], c[1171]);
HA HA_82(r[812], r[813], r[1172], c[1172]);
FA FA_1090(c[598], r[599], r[600], r[1173], c[1173]);
FA FA_1091(r[601], c[812], c[813], r[1174], c[1174]);
HA HA_83(c[814], r[815], r[1175], c[1175]);
FA FA_1092(c[601], r[602], r[603], r[1176], c[1176]);
FA FA_1093(r[604], c[815], c[816], r[1177], c[1177]);
HA HA_84(c[817], r[818], r[1178], c[1178]);
FA FA_1094(c[604], r[605], r[606], r[1179], c[1179]);
FA FA_1095(r[607], c[818], c[819], r[1180], c[1180]);
HA HA_85(c[820], r[821], r[1181], c[1181]);
FA FA_1096(c[607], r[608], r[609], r[1182], c[1182]);
FA FA_1097(r[610], c[821], c[822], r[1183], c[1183]);
FA FA_1098(c[610], r[611], r[612], r[1184], c[1184]);
FA FA_1099(r[613], c[824], c[825], r[1185], c[1185]);
FA FA_1100(c[613], r[614], r[615], r[1186], c[1186]);
FA FA_1101(r[616], c[827], c[828], r[1187], c[1187]);
FA FA_1102(r[617], r[618], r[619], r[1188], c[1188]);
FA FA_1103(r[620], c[830], c[831], r[1189], c[1189]);
FA FA_1104(r[621], r[622], r[623], r[1190], c[1190]);
FA FA_1105(r[624], c[833], c[834], r[1191], c[1191]);
FA FA_1106(c[622], c[623], c[624], r[1192], c[1192]);
FA FA_1107(r[625], r[626], r[627], r[1193], c[1193]);
FA FA_1108(r[628], c[836], c[837], r[1194], c[1194]);
FA FA_1109(c[626], c[627], c[628], r[1195], c[1195]);
FA FA_1110(r[629], r[630], r[631], r[1196], c[1196]);
FA FA_1111(r[632], c[839], c[840], r[1197], c[1197]);
FA FA_1112(c[630], c[631], c[632], r[1198], c[1198]);
FA FA_1113(r[633], r[634], r[635], r[1199], c[1199]);
FA FA_1114(r[636], c[842], c[843], r[1200], c[1200]);
FA FA_1115(c[635], c[636], r[637], r[1201], c[1201]);
FA FA_1116(r[638], r[639], r[640], r[1202], c[1202]);
FA FA_1117(c[845], c[846], c[847], r[1203], c[1203]);
FA FA_1118(c[640], r[641], r[642], r[1204], c[1204]);
FA FA_1119(r[643], r[644], c[848], r[1205], c[1205]);
FA FA_1120(c[849], c[850], c[851], r[1206], c[1206]);
FA FA_1121(r[646], r[647], r[648], r[1207], c[1207]);
FA FA_1122(c[852], c[853], c[854], r[1208], c[1208]);
FA FA_1123(c[855], r[856], r[857], r[1209], c[1209]);
FA FA_1124(c[648], r[649], r[650], r[1210], c[1210]);
FA FA_1125(r[651], r[652], c[856], r[1211], c[1211]);
FA FA_1126(c[857], c[858], c[859], r[1212], c[1212]);
FA FA_1127(c[652], r[653], r[654], r[1213], c[1213]);
FA FA_1128(r[655], r[656], c[861], r[1214], c[1214]);
FA FA_1129(c[862], c[863], c[864], r[1215], c[1215]);
FA FA_1130(c[656], r[657], r[658], r[1216], c[1216]);
FA FA_1131(r[659], r[660], r[661], r[1217], c[1217]);
FA FA_1132(c[865], c[866], c[867], r[1218], c[1218]);
FA FA_1133(c[661], r[662], r[663], r[1219], c[1219]);
FA FA_1134(r[664], r[665], r[666], r[1220], c[1220]);
FA FA_1135(c[870], c[871], c[872], r[1221], c[1221]);
FA FA_1136(c[666], r[667], r[668], r[1222], c[1222]);
FA FA_1137(r[669], r[670], r[671], r[1223], c[1223]);
FA FA_1138(c[874], c[875], c[876], r[1224], c[1224]);
FA FA_1139(r[672], r[673], r[674], r[1225], c[1225]);
FA FA_1140(r[675], r[676], r[677], r[1226], c[1226]);
FA FA_1141(c[878], c[879], c[880], r[1227], c[1227]);
FA FA_1142(c[674], c[675], c[676], r[1228], c[1228]);
FA FA_1143(c[677], r[678], r[679], r[1229], c[1229]);
FA FA_1144(r[680], r[681], r[682], r[1230], c[1230]);
FA FA_1145(c[682], r[683], r[684], r[1231], c[1231]);
FA FA_1146(r[685], r[686], r[687], r[1232], c[1232]);
FA FA_1147(c[886], c[887], c[888], r[1233], c[1233]);
HA HA_86(c[889], r[890], r[1234], c[1234]);
FA FA_1148(c[685], c[686], c[687], r[1235], c[1235]);
FA FA_1149(r[688], r[689], r[690], r[1236], c[1236]);
FA FA_1150(r[691], r[692], c[890], r[1237], c[1237]);
HA HA_87(c[891], c[892], r[1238], c[1238]);
FA FA_1151(c[690], c[691], c[692], r[1239], c[1239]);
FA FA_1152(r[693], r[694], r[695], r[1240], c[1240]);
FA FA_1153(r[696], r[697], r[698], r[1241], c[1241]);
HA HA_88(c[894], c[895], r[1242], c[1242]);
FA FA_1154(c[695], c[696], c[697], r[1243], c[1243]);
FA FA_1155(c[698], r[699], r[700], r[1244], c[1244]);
FA FA_1156(r[701], r[702], r[703], r[1245], c[1245]);
FA FA_1157(c[898], c[899], c[900], r[1246], c[1246]);
FA FA_1158(c[703], r[704], r[705], r[1247], c[1247]);
FA FA_1159(r[706], r[707], r[708], r[1248], c[1248]);
FA FA_1160(r[709], c[902], c[903], r[1249], c[1249]);
FA FA_1161(c[904], c[905], c[906], r[1250], c[1250]);
FA FA_1162(c[706], c[707], c[708], r[1251], c[1251]);
FA FA_1163(c[709], r[710], r[711], r[1252], c[1252]);
FA FA_1164(r[712], r[713], r[714], r[1253], c[1253]);
FA FA_1165(c[907], c[908], c[909], r[1254], c[1254]);
HA HA_89(c[910], c[911], r[1255], c[1255]);
FA FA_1166(c[714], r[715], r[716], r[1256], c[1256]);
FA FA_1167(r[717], r[718], r[719], r[1257], c[1257]);
FA FA_1168(r[720], c[913], c[914], r[1258], c[1258]);
FA FA_1169(c[915], c[916], c[917], r[1259], c[1259]);
FA FA_1170(c[717], c[718], c[719], r[1260], c[1260]);
FA FA_1171(c[720], r[721], r[722], r[1261], c[1261]);
FA FA_1172(r[723], r[724], r[725], r[1262], c[1262]);
FA FA_1173(r[726], c[918], c[919], r[1263], c[1263]);
FA FA_1174(c[723], c[724], c[725], r[1264], c[1264]);
FA FA_1175(c[726], r[727], r[728], r[1265], c[1265]);
FA FA_1176(r[729], r[730], r[731], r[1266], c[1266]);
FA FA_1177(r[732], c[924], c[925], r[1267], c[1267]);
HA HA_90(c[926], c[927], r[1268], c[1268]);
FA FA_1178(c[730], c[731], c[732], r[1269], c[1269]);
FA FA_1179(r[733], r[734], r[735], r[1270], c[1270]);
FA FA_1180(r[736], r[737], r[738], r[1271], c[1271]);
FA FA_1181(r[739], c[929], c[930], r[1272], c[1272]);
FA FA_1182(c[736], c[737], c[738], r[1273], c[1273]);
FA FA_1183(c[739], r[740], r[741], r[1274], c[1274]);
FA FA_1184(r[742], r[743], r[744], r[1275], c[1275]);
FA FA_1185(r[745], c[934], c[935], r[1276], c[1276]);
FA FA_1186(c[743], c[744], c[745], r[1277], c[1277]);
FA FA_1187(r[746], r[747], r[748], r[1278], c[1278]);
FA FA_1188(r[749], r[750], r[751], r[1279], c[1279]);
FA FA_1189(r[752], c[939], c[940], r[1280], c[1280]);
FA FA_1190(c[751], c[752], r[753], r[1281], c[1281]);
FA FA_1191(r[754], r[755], r[756], r[1282], c[1282]);
FA FA_1192(r[757], r[758], c[945], r[1283], c[1283]);
FA FA_1193(c[946], c[947], c[948], r[1284], c[1284]);
FA FA_1194(c[756], c[757], c[758], r[1285], c[1285]);
FA FA_1195(r[759], r[760], r[761], r[1286], c[1286]);
FA FA_1196(r[762], r[763], r[764], r[1287], c[1287]);
FA FA_1197(r[765], c[950], c[951], r[1288], c[1288]);
FA FA_1198(c[765], r[766], r[767], r[1289], c[1289]);
FA FA_1199(r[768], r[769], r[770], r[1290], c[1290]);
FA FA_1200(r[771], r[772], c[956], r[1291], c[1291]);
FA FA_1201(c[957], c[958], c[959], r[1292], c[1292]);
HA HA_91(r[968], r[1139], r[1293], c[1293]);
FA FA_1202(r[1140], r[1141], c[1293], r[1294], c[1294]);
FA FA_1203(r[970], c[1140], c[1141], r[1295], c[1295]);
HA HA_92(r[1142], c[1294], r[1296], c[1296]);
FA FA_1204(r[971], r[972], c[1142], r[1297], c[1297]);
FA FA_1205(c[972], r[973], c[1143], r[1298], c[1298]);
HA HA_93(r[1144], c[1297], r[1299], c[1299]);
FA FA_1206(c[973], r[974], c[1144], r[1300], c[1300]);
FA FA_1207(r[975], r[976], c[1145], r[1301], c[1301]);
FA FA_1208(c[976], r[977], c[1147], r[1302], c[1302]);
FA FA_1209(c[786], r[787], c[977], r[1303], c[1303]);
HA HA_94(r[978], c[1148], r[1304], c[1304]);
FA FA_1210(c[787], r[788], r[789], r[1305], c[1305]);
FA FA_1211(c[789], r[790], r[791], r[1306], c[1306]);
HA HA_95(c[979], r[980], r[1307], c[1307]);
FA FA_1212(r[792], r[793], r[794], r[1308], c[1308]);
FA FA_1213(r[795], r[796], c[981], r[1309], c[1309]);
HA HA_96(r[982], r[983], r[1310], c[1310]);
FA FA_1214(r[798], c[982], c[983], r[1311], c[1311]);
FA FA_1215(c[984], c[985], c[986], r[1312], c[1312]);
FA FA_1216(c[988], r[989], r[990], r[1313], c[1313]);
FA FA_1217(c[989], c[990], c[991], r[1314], c[1314]);
FA FA_1218(c[993], r[994], r[995], r[1315], c[1315]);
FA FA_1219(c[994], c[995], c[996], r[1316], c[1316]);
FA FA_1220(r[997], r[998], r[999], r[1317], c[1317]);
FA FA_1221(c[999], r[1000], r[1001], r[1318], c[1318]);
HA HA_97(r[1002], c[1165], r[1319], c[1319]);
FA FA_1222(r[814], c[1000], c[1001], r[1320], c[1320]);
FA FA_1223(c[1002], r[1003], r[1004], r[1321], c[1321]);
HA HA_98(c[1167], c[1168], r[1322], c[1322]);
FA FA_1224(r[816], r[817], c[1003], r[1323], c[1323]);
FA FA_1225(c[1004], r[1005], r[1006], r[1324], c[1324]);
FA FA_1226(r[819], r[820], c[1005], r[1325], c[1325]);
FA FA_1227(c[1006], r[1007], r[1008], r[1326], c[1326]);
HA HA_99(c[1173], c[1174], r[1327], c[1327]);
FA FA_1228(r[822], r[823], c[1007], r[1328], c[1328]);
FA FA_1229(c[1008], r[1009], r[1010], r[1329], c[1329]);
FA FA_1230(c[823], r[824], r[825], r[1330], c[1330]);
FA FA_1231(r[826], c[1009], c[1010], r[1331], c[1331]);
FA FA_1232(c[826], r[827], r[828], r[1332], c[1332]);
FA FA_1233(r[829], c[1011], c[1012], r[1333], c[1333]);
FA FA_1234(c[829], r[830], r[831], r[1334], c[1334]);
FA FA_1235(r[832], c[1014], c[1015], r[1335], c[1335]);
FA FA_1236(c[832], r[833], r[834], r[1336], c[1336]);
FA FA_1237(r[835], c[1017], c[1018], r[1337], c[1337]);
FA FA_1238(c[835], r[836], r[837], r[1338], c[1338]);
FA FA_1239(r[838], c[1020], c[1021], r[1339], c[1339]);
FA FA_1240(c[838], r[839], r[840], r[1340], c[1340]);
FA FA_1241(r[841], c[1023], c[1024], r[1341], c[1341]);
HA HA_100(c[1025], r[1026], r[1342], c[1342]);
FA FA_1242(c[841], r[842], r[843], r[1343], c[1343]);
FA FA_1243(r[844], c[1026], c[1027], r[1344], c[1344]);
FA FA_1244(c[844], r[845], r[846], r[1345], c[1345]);
FA FA_1245(r[847], c[1029], c[1030], r[1346], c[1346]);
FA FA_1246(r[848], r[849], r[850], r[1347], c[1347]);
FA FA_1247(r[851], c[1032], c[1033], r[1348], c[1348]);
FA FA_1248(r[852], r[853], r[854], r[1349], c[1349]);
FA FA_1249(r[855], c[1035], c[1036], r[1350], c[1350]);
FA FA_1250(r[858], r[859], r[860], r[1351], c[1351]);
FA FA_1251(c[1038], c[1039], c[1040], r[1352], c[1352]);
FA FA_1252(c[860], r[861], r[862], r[1353], c[1353]);
FA FA_1253(r[863], r[864], c[1041], r[1354], c[1354]);
FA FA_1254(c[1042], c[1043], c[1044], r[1355], c[1355]);
FA FA_1255(r[865], r[866], r[867], r[1356], c[1356]);
FA FA_1256(r[868], r[869], c[1045], r[1357], c[1357]);
FA FA_1257(c[1046], c[1047], c[1048], r[1358], c[1358]);
FA FA_1258(c[868], c[869], r[870], r[1359], c[1359]);
FA FA_1259(r[871], r[872], r[873], r[1360], c[1360]);
FA FA_1260(c[1049], c[1050], c[1051], r[1361], c[1361]);
FA FA_1261(c[873], r[874], r[875], r[1362], c[1362]);
FA FA_1262(r[876], r[877], c[1052], r[1363], c[1363]);
FA FA_1263(c[1053], c[1054], c[1055], r[1364], c[1364]);
FA FA_1264(c[877], r[878], r[879], r[1365], c[1365]);
FA FA_1265(r[880], r[881], c[1056], r[1366], c[1366]);
FA FA_1266(c[1057], c[1058], c[1059], r[1367], c[1367]);
FA FA_1267(c[881], r[882], r[883], r[1368], c[1368]);
FA FA_1268(r[884], r[885], c[1060], r[1369], c[1369]);
FA FA_1269(c[1061], c[1062], c[1063], r[1370], c[1370]);
FA FA_1270(c[882], c[883], c[884], r[1371], c[1371]);
FA FA_1271(c[885], r[886], r[887], r[1372], c[1372]);
FA FA_1272(r[888], r[889], c[1064], r[1373], c[1373]);
FA FA_1273(r[891], r[892], r[893], r[1374], c[1374]);
FA FA_1274(c[1068], c[1069], c[1070], r[1375], c[1375]);
FA FA_1275(c[1071], r[1072], r[1073], r[1376], c[1376]);
FA FA_1276(c[893], r[894], r[895], r[1377], c[1377]);
FA FA_1277(r[896], r[897], c[1072], r[1378], c[1378]);
FA FA_1278(c[1073], c[1074], c[1075], r[1379], c[1379]);
FA FA_1279(c[896], c[897], r[898], r[1380], c[1380]);
FA FA_1280(r[899], r[900], r[901], r[1381], c[1381]);
FA FA_1281(c[1077], c[1078], c[1079], r[1382], c[1382]);
FA FA_1282(c[901], r[902], r[903], r[1383], c[1383]);
FA FA_1283(r[904], r[905], r[906], r[1384], c[1384]);
FA FA_1284(c[1081], c[1082], c[1083], r[1385], c[1385]);
FA FA_1285(r[907], r[908], r[909], r[1386], c[1386]);
FA FA_1286(r[910], r[911], r[912], r[1387], c[1387]);
FA FA_1287(c[1085], c[1086], c[1087], r[1388], c[1388]);
FA FA_1288(c[912], r[913], r[914], r[1389], c[1389]);
FA FA_1289(r[915], r[916], r[917], r[1390], c[1390]);
FA FA_1290(c[1089], c[1090], c[1091], r[1391], c[1391]);
HA HA_101(c[1092], r[1093], r[1392], c[1392]);
FA FA_1291(r[918], r[919], r[920], r[1393], c[1393]);
FA FA_1292(r[921], r[922], r[923], r[1394], c[1394]);
FA FA_1293(c[1093], c[1094], c[1095], r[1395], c[1395]);
FA FA_1294(c[920], c[921], c[922], r[1396], c[1396]);
FA FA_1295(c[923], r[924], r[925], r[1397], c[1397]);
FA FA_1296(r[926], r[927], r[928], r[1398], c[1398]);
FA FA_1297(c[928], r[929], r[930], r[1399], c[1399]);
FA FA_1298(r[931], r[932], r[933], r[1400], c[1400]);
FA FA_1299(c[1101], c[1102], c[1103], r[1401], c[1401]);
HA HA_102(c[1104], r[1105], r[1402], c[1402]);
FA FA_1300(c[931], c[932], c[933], r[1403], c[1403]);
FA FA_1301(r[934], r[935], r[936], r[1404], c[1404]);
FA FA_1302(r[937], r[938], c[1105], r[1405], c[1405]);
HA HA_103(c[1106], c[1107], r[1406], c[1406]);
FA FA_1303(c[936], c[937], c[938], r[1407], c[1407]);
FA FA_1304(r[939], r[940], r[941], r[1408], c[1408]);
FA FA_1305(r[942], r[943], r[944], r[1409], c[1409]);
HA HA_104(c[1109], c[1110], r[1410], c[1410]);
FA FA_1306(c[941], c[942], c[943], r[1411], c[1411]);
FA FA_1307(c[944], r[945], r[946], r[1412], c[1412]);
FA FA_1308(r[947], r[948], r[949], r[1413], c[1413]);
FA FA_1309(c[1113], c[1114], c[1115], r[1414], c[1414]);
FA FA_1310(c[949], r[950], r[951], r[1415], c[1415]);
FA FA_1311(r[952], r[953], r[954], r[1416], c[1416]);
FA FA_1312(r[955], c[1117], c[1118], r[1417], c[1417]);
FA FA_1313(c[1119], c[1120], c[1121], r[1418], c[1418]);
FA FA_1314(c[952], c[953], c[954], r[1419], c[1419]);
FA FA_1315(c[955], r[956], r[957], r[1420], c[1420]);
FA FA_1316(r[958], r[959], r[960], r[1421], c[1421]);
FA FA_1317(c[1122], c[1123], c[1124], r[1422], c[1422]);
HA HA_105(c[1125], c[1126], r[1423], c[1423]);
FA FA_1318(c[960], r[961], r[962], r[1424], c[1424]);
FA FA_1319(r[963], r[964], r[965], r[1425], c[1425]);
FA FA_1320(r[966], c[1128], c[1129], r[1426], c[1426]);
FA FA_1321(c[1130], c[1131], c[1132], r[1427], c[1427]);
HA HA_106(r[1295], r[1296], r[1428], c[1428]);
FA FA_1322(r[1143], c[1295], c[1296], r[1429], c[1429]);
HA HA_107(r[1297], c[1428], r[1430], c[1430]);
FA FA_1323(r[1298], r[1299], c[1429], r[1431], c[1431]);
FA FA_1324(r[1145], r[1146], c[1298], r[1432], c[1432]);
FA FA_1325(c[1146], r[1147], c[1300], r[1433], c[1433]);
HA HA_108(r[1301], c[1432], r[1434], c[1434]);
FA FA_1326(r[1148], r[1149], c[1301], r[1435], c[1435]);
FA FA_1327(c[1149], r[1150], c[1302], r[1436], c[1436]);
FA FA_1328(c[978], r[979], c[1150], r[1437], c[1437]);
HA HA_109(r[1151], c[1303], r[1438], c[1438]);
FA FA_1329(c[1151], r[1152], c[1305], r[1439], c[1439]);
FA FA_1330(c[980], r[981], c[1152], r[1440], c[1440]);
HA HA_110(r[1153], c[1306], r[1441], c[1441]);
FA FA_1331(c[1153], r[1154], c[1308], r[1442], c[1442]);
FA FA_1332(r[984], r[985], r[986], r[1443], c[1443]);
FA FA_1333(r[987], r[988], c[1155], r[1444], c[1444]);
HA HA_111(r[1156], r[1157], r[1445], c[1445]);
FA FA_1334(r[991], c[1156], c[1157], r[1446], c[1446]);
FA FA_1335(r[992], r[993], c[1158], r[1447], c[1447]);
FA FA_1336(r[996], c[1160], c[1161], r[1448], c[1448]);
FA FA_1337(c[1162], c[1163], c[1164], r[1449], c[1449]);
FA FA_1338(c[1166], r[1167], r[1168], r[1450], c[1450]);
FA FA_1339(c[1169], r[1170], r[1171], r[1451], c[1451]);
FA FA_1340(c[1170], c[1171], c[1172], r[1452], c[1452]);
FA FA_1341(r[1173], r[1174], r[1175], r[1453], c[1453]);
FA FA_1342(c[1175], r[1176], r[1177], r[1454], c[1454]);
HA HA_112(r[1178], c[1323], r[1455], c[1455]);
FA FA_1343(c[1176], c[1177], c[1178], r[1456], c[1456]);
FA FA_1344(r[1179], r[1180], r[1181], r[1457], c[1457]);
FA FA_1345(r[1011], r[1012], r[1013], r[1458], c[1458]);
FA FA_1346(c[1179], c[1180], c[1181], r[1459], c[1459]);
HA HA_113(r[1182], r[1183], r[1460], c[1460]);
FA FA_1347(c[1013], r[1014], r[1015], r[1461], c[1461]);
FA FA_1348(r[1016], c[1182], c[1183], r[1462], c[1462]);
FA FA_1349(c[1016], r[1017], r[1018], r[1463], c[1463]);
FA FA_1350(r[1019], c[1184], c[1185], r[1464], c[1464]);
HA HA_114(r[1186], r[1187], r[1465], c[1465]);
FA FA_1351(c[1019], r[1020], r[1021], r[1466], c[1466]);
FA FA_1352(r[1022], c[1186], c[1187], r[1467], c[1467]);
FA FA_1353(c[1022], r[1023], r[1024], r[1468], c[1468]);
FA FA_1354(r[1025], c[1188], c[1189], r[1469], c[1469]);
HA HA_115(r[1190], r[1191], r[1470], c[1470]);
FA FA_1355(r[1027], r[1028], c[1190], r[1471], c[1471]);
FA FA_1356(c[1191], r[1192], r[1193], r[1472], c[1472]);
FA FA_1357(c[1028], r[1029], r[1030], r[1473], c[1473]);
FA FA_1358(r[1031], c[1192], c[1193], r[1474], c[1474]);
HA HA_116(c[1194], r[1195], r[1475], c[1475]);
FA FA_1359(c[1031], r[1032], r[1033], r[1476], c[1476]);
FA FA_1360(r[1034], c[1195], c[1196], r[1477], c[1477]);
HA HA_117(c[1197], r[1198], r[1478], c[1478]);
FA FA_1361(c[1034], r[1035], r[1036], r[1479], c[1479]);
FA FA_1362(r[1037], c[1198], c[1199], r[1480], c[1480]);
HA HA_118(c[1200], r[1201], r[1481], c[1481]);
FA FA_1363(c[1037], r[1038], r[1039], r[1482], c[1482]);
FA FA_1364(r[1040], c[1201], c[1202], r[1483], c[1483]);
HA HA_119(c[1203], r[1204], r[1484], c[1484]);
FA FA_1365(r[1041], r[1042], r[1043], r[1485], c[1485]);
FA FA_1366(r[1044], c[1204], c[1205], r[1486], c[1486]);
HA HA_120(c[1206], r[1207], r[1487], c[1487]);
FA FA_1367(r[1045], r[1046], r[1047], r[1488], c[1488]);
FA FA_1368(r[1048], c[1207], c[1208], r[1489], c[1489]);
FA FA_1369(r[1049], r[1050], r[1051], r[1490], c[1490]);
FA FA_1370(c[1210], c[1211], c[1212], r[1491], c[1491]);
HA HA_121(r[1213], r[1214], r[1492], c[1492]);
FA FA_1371(r[1052], r[1053], r[1054], r[1493], c[1493]);
FA FA_1372(r[1055], c[1213], c[1214], r[1494], c[1494]);
FA FA_1373(r[1056], r[1057], r[1058], r[1495], c[1495]);
FA FA_1374(r[1059], c[1216], c[1217], r[1496], c[1496]);
FA FA_1375(r[1060], r[1061], r[1062], r[1497], c[1497]);
FA FA_1376(r[1063], c[1219], c[1220], r[1498], c[1498]);
FA FA_1377(r[1064], r[1065], r[1066], r[1499], c[1499]);
FA FA_1378(r[1067], c[1222], c[1223], r[1500], c[1500]);
FA FA_1379(c[1065], c[1066], c[1067], r[1501], c[1501]);
FA FA_1380(r[1068], r[1069], r[1070], r[1502], c[1502]);
FA FA_1381(r[1071], c[1225], c[1226], r[1503], c[1503]);
FA FA_1382(r[1074], r[1075], r[1076], r[1504], c[1504]);
FA FA_1383(c[1228], c[1229], c[1230], r[1505], c[1505]);
FA FA_1384(c[1076], r[1077], r[1078], r[1506], c[1506]);
FA FA_1385(r[1079], r[1080], c[1231], r[1507], c[1507]);
FA FA_1386(c[1232], c[1233], c[1234], r[1508], c[1508]);
FA FA_1387(c[1080], r[1081], r[1082], r[1509], c[1509]);
FA FA_1388(r[1083], r[1084], c[1235], r[1510], c[1510]);
FA FA_1389(c[1236], c[1237], c[1238], r[1511], c[1511]);
FA FA_1390(c[1084], r[1085], r[1086], r[1512], c[1512]);
FA FA_1391(r[1087], r[1088], c[1239], r[1513], c[1513]);
FA FA_1392(c[1240], c[1241], c[1242], r[1514], c[1514]);
FA FA_1393(c[1088], r[1089], r[1090], r[1515], c[1515]);
FA FA_1394(r[1091], r[1092], c[1243], r[1516], c[1516]);
FA FA_1395(c[1244], c[1245], c[1246], r[1517], c[1517]);
FA FA_1396(r[1094], r[1095], r[1096], r[1518], c[1518]);
FA FA_1397(c[1247], c[1248], c[1249], r[1519], c[1519]);
FA FA_1398(c[1250], r[1251], r[1252], r[1520], c[1520]);
FA FA_1399(c[1096], r[1097], r[1098], r[1521], c[1521]);
FA FA_1400(r[1099], r[1100], c[1251], r[1522], c[1522]);
FA FA_1401(c[1252], c[1253], c[1254], r[1523], c[1523]);
FA FA_1402(c[1097], c[1098], c[1099], r[1524], c[1524]);
FA FA_1403(c[1100], r[1101], r[1102], r[1525], c[1525]);
FA FA_1404(r[1103], r[1104], c[1256], r[1526], c[1526]);
FA FA_1405(r[1106], r[1107], r[1108], r[1527], c[1527]);
FA FA_1406(c[1260], c[1261], c[1262], r[1528], c[1528]);
FA FA_1407(c[1263], r[1264], r[1265], r[1529], c[1529]);
FA FA_1408(c[1108], r[1109], r[1110], r[1530], c[1530]);
FA FA_1409(r[1111], r[1112], c[1264], r[1531], c[1531]);
FA FA_1410(c[1265], c[1266], c[1267], r[1532], c[1532]);
FA FA_1411(c[1111], c[1112], r[1113], r[1533], c[1533]);
FA FA_1412(r[1114], r[1115], r[1116], r[1534], c[1534]);
FA FA_1413(c[1269], c[1270], c[1271], r[1535], c[1535]);
FA FA_1414(c[1116], r[1117], r[1118], r[1536], c[1536]);
FA FA_1415(r[1119], r[1120], r[1121], r[1537], c[1537]);
FA FA_1416(c[1273], c[1274], c[1275], r[1538], c[1538]);
FA FA_1417(r[1122], r[1123], r[1124], r[1539], c[1539]);
FA FA_1418(r[1125], r[1126], r[1127], r[1540], c[1540]);
FA FA_1419(c[1277], c[1278], c[1279], r[1541], c[1541]);
FA FA_1420(c[1127], r[1128], r[1129], r[1542], c[1542]);
FA FA_1421(r[1130], r[1131], r[1132], r[1543], c[1543]);
FA FA_1422(c[1281], c[1282], c[1283], r[1544], c[1544]);
HA HA_122(c[1284], r[1285], r[1545], c[1545]);
FA FA_1423(r[1133], r[1134], r[1135], r[1546], c[1546]);
FA FA_1424(r[1136], r[1137], r[1138], r[1547], c[1547]);
FA FA_1425(c[1285], c[1286], c[1287], r[1548], c[1548]);
HA HA_123(r[1429], r[1430], r[1549], c[1549]);
FA FA_1426(c[1430], r[1431], c[1549], r[1550], c[1550]);
FA FA_1427(c[1299], r[1300], c[1431], r[1551], c[1551]);
HA HA_124(r[1432], c[1550], r[1552], c[1552]);
FA FA_1428(r[1433], r[1434], c[1551], r[1553], c[1553]);
FA FA_1429(r[1302], c[1433], c[1434], r[1554], c[1554]);
HA HA_125(r[1435], c[1553], r[1555], c[1555]);
FA FA_1430(r[1303], r[1304], c[1435], r[1556], c[1556]);
FA FA_1431(c[1304], r[1305], c[1436], r[1557], c[1557]);
FA FA_1432(r[1306], r[1307], c[1437], r[1558], c[1558]);
FA FA_1433(c[1307], r[1308], c[1439], r[1559], c[1559]);
FA FA_1434(r[1309], r[1310], c[1440], r[1560], c[1560]);
FA FA_1435(c[1154], r[1155], c[1309], r[1561], c[1561]);
HA HA_126(c[1310], r[1311], r[1562], c[1562]);
FA FA_1436(c[1311], r[1312], c[1443], r[1563], c[1563]);
FA FA_1437(r[1158], r[1159], c[1312], r[1564], c[1564]);
HA HA_127(r[1313], c[1444], r[1565], c[1565]);
FA FA_1438(c[1159], r[1160], r[1161], r[1566], c[1566]);
FA FA_1439(r[1162], r[1163], r[1164], r[1567], c[1567]);
HA HA_128(c[1314], r[1315], r[1568], c[1568]);
FA FA_1440(r[1165], r[1166], c[1315], r[1569], c[1569]);
FA FA_1441(r[1169], c[1316], c[1317], r[1570], c[1570]);
HA HA_129(r[1318], r[1319], r[1571], c[1571]);
FA FA_1442(r[1172], c[1318], c[1319], r[1572], c[1572]);
FA FA_1443(c[1320], c[1321], c[1322], r[1573], c[1573]);
FA FA_1444(c[1324], r[1325], r[1326], r[1574], c[1574]);
FA FA_1445(c[1325], c[1326], c[1327], r[1575], c[1575]);
FA FA_1446(c[1328], c[1329], r[1330], r[1576], c[1576]);
FA FA_1447(r[1184], r[1185], c[1330], r[1577], c[1577]);
FA FA_1448(c[1331], r[1332], r[1333], r[1578], c[1578]);
FA FA_1449(c[1332], c[1333], r[1334], r[1579], c[1579]);
HA HA_130(r[1335], c[1461], r[1580], c[1580]);
FA FA_1450(r[1188], r[1189], c[1334], r[1581], c[1581]);
FA FA_1451(c[1335], r[1336], r[1337], r[1582], c[1582]);
FA FA_1452(c[1336], c[1337], r[1338], r[1583], c[1583]);
HA HA_131(r[1339], c[1466], r[1584], c[1584]);
FA FA_1453(r[1194], c[1338], c[1339], r[1585], c[1585]);
FA FA_1454(r[1340], r[1341], r[1342], r[1586], c[1586]);
FA FA_1455(r[1196], r[1197], c[1340], r[1587], c[1587]);
FA FA_1456(c[1341], c[1342], r[1343], r[1588], c[1588]);
HA HA_132(r[1344], c[1471], r[1589], c[1589]);
FA FA_1457(r[1199], r[1200], c[1343], r[1590], c[1590]);
FA FA_1458(c[1344], r[1345], r[1346], r[1591], c[1591]);
FA FA_1459(r[1202], r[1203], c[1345], r[1592], c[1592]);
FA FA_1460(c[1346], r[1347], r[1348], r[1593], c[1593]);
HA HA_133(c[1476], c[1477], r[1594], c[1594]);
FA FA_1461(r[1205], r[1206], c[1347], r[1595], c[1595]);
FA FA_1462(c[1348], r[1349], r[1350], r[1596], c[1596]);
FA FA_1463(r[1208], r[1209], c[1349], r[1597], c[1597]);
FA FA_1464(c[1350], r[1351], r[1352], r[1598], c[1598]);
HA HA_134(c[1482], c[1483], r[1599], c[1599]);
FA FA_1465(c[1209], r[1210], r[1211], r[1600], c[1600]);
FA FA_1466(r[1212], c[1351], c[1352], r[1601], c[1601]);
HA HA_135(r[1353], r[1354], r[1602], c[1602]);
FA FA_1467(r[1215], c[1353], c[1354], r[1603], c[1603]);
FA FA_1468(c[1355], r[1356], r[1357], r[1604], c[1604]);
FA FA_1469(c[1215], r[1216], r[1217], r[1605], c[1605]);
FA FA_1470(r[1218], c[1356], c[1357], r[1606], c[1606]);
HA HA_136(c[1358], r[1359], r[1607], c[1607]);
FA FA_1471(c[1218], r[1219], r[1220], r[1608], c[1608]);
FA FA_1472(r[1221], c[1359], c[1360], r[1609], c[1609]);
HA HA_137(c[1361], r[1362], r[1610], c[1610]);
FA FA_1473(c[1221], r[1222], r[1223], r[1611], c[1611]);
FA FA_1474(r[1224], c[1362], c[1363], r[1612], c[1612]);
HA HA_138(c[1364], r[1365], r[1613], c[1613]);
FA FA_1475(c[1224], r[1225], r[1226], r[1614], c[1614]);
FA FA_1476(r[1227], c[1365], c[1366], r[1615], c[1615]);
HA HA_139(c[1367], r[1368], r[1616], c[1616]);
FA FA_1477(c[1227], r[1228], r[1229], r[1617], c[1617]);
FA FA_1478(r[1230], c[1368], c[1369], r[1618], c[1618]);
FA FA_1479(r[1231], r[1232], r[1233], r[1619], c[1619]);
FA FA_1480(r[1234], c[1371], c[1372], r[1620], c[1620]);
HA HA_140(c[1373], r[1374], r[1621], c[1621]);
FA FA_1481(r[1235], r[1236], r[1237], r[1622], c[1622]);
FA FA_1482(r[1238], c[1374], c[1375], r[1623], c[1623]);
FA FA_1483(r[1239], r[1240], r[1241], r[1624], c[1624]);
FA FA_1484(r[1242], c[1377], c[1378], r[1625], c[1625]);
FA FA_1485(r[1243], r[1244], r[1245], r[1626], c[1626]);
FA FA_1486(r[1246], c[1380], c[1381], r[1627], c[1627]);
FA FA_1487(r[1247], r[1248], r[1249], r[1628], c[1628]);
FA FA_1488(r[1250], c[1383], c[1384], r[1629], c[1629]);
FA FA_1489(r[1253], r[1254], r[1255], r[1630], c[1630]);
FA FA_1490(c[1386], c[1387], c[1388], r[1631], c[1631]);
FA FA_1491(c[1255], r[1256], r[1257], r[1632], c[1632]);
FA FA_1492(r[1258], r[1259], c[1389], r[1633], c[1633]);
HA HA_141(c[1390], c[1391], r[1634], c[1634]);
FA FA_1493(c[1257], c[1258], c[1259], r[1635], c[1635]);
FA FA_1494(r[1260], r[1261], r[1262], r[1636], c[1636]);
FA FA_1495(r[1263], c[1393], c[1394], r[1637], c[1637]);
FA FA_1496(r[1266], r[1267], r[1268], r[1638], c[1638]);
FA FA_1497(c[1396], c[1397], c[1398], r[1639], c[1639]);
FA FA_1498(c[1268], r[1269], r[1270], r[1640], c[1640]);
FA FA_1499(r[1271], r[1272], c[1399], r[1641], c[1641]);
FA FA_1500(c[1400], c[1401], c[1402], r[1642], c[1642]);
FA FA_1501(c[1272], r[1273], r[1274], r[1643], c[1643]);
FA FA_1502(r[1275], r[1276], c[1403], r[1644], c[1644]);
FA FA_1503(c[1404], c[1405], c[1406], r[1645], c[1645]);
FA FA_1504(c[1276], r[1277], r[1278], r[1646], c[1646]);
FA FA_1505(r[1279], r[1280], c[1407], r[1647], c[1647]);
FA FA_1506(c[1408], c[1409], c[1410], r[1648], c[1648]);
FA FA_1507(c[1280], r[1281], r[1282], r[1649], c[1649]);
FA FA_1508(r[1283], r[1284], c[1411], r[1650], c[1650]);
FA FA_1509(c[1412], c[1413], c[1414], r[1651], c[1651]);
FA FA_1510(r[1286], r[1287], r[1288], r[1652], c[1652]);
FA FA_1511(c[1415], c[1416], c[1417], r[1653], c[1653]);
FA FA_1512(c[1418], r[1419], r[1420], r[1654], c[1654]);
FA FA_1513(c[1288], r[1289], r[1290], r[1655], c[1655]);
FA FA_1514(r[1291], r[1292], c[1419], r[1656], c[1656]);
FA FA_1515(c[1420], c[1421], c[1422], r[1657], c[1657]);
HA HA_142(r[1551], r[1552], r[1658], c[1658]);
FA FA_1516(c[1552], r[1553], c[1658], r[1659], c[1659]);
FA FA_1517(r[1554], r[1555], c[1659], r[1660], c[1660]);
FA FA_1518(r[1436], c[1554], c[1555], r[1661], c[1661]);
HA HA_143(r[1556], c[1660], r[1662], c[1662]);
FA FA_1519(r[1437], r[1438], c[1556], r[1663], c[1663]);
FA FA_1520(c[1438], r[1439], c[1557], r[1664], c[1664]);
HA HA_144(r[1558], c[1663], r[1665], c[1665]);
FA FA_1521(r[1440], r[1441], c[1558], r[1666], c[1666]);
FA FA_1522(c[1441], r[1442], c[1559], r[1667], c[1667]);
HA HA_145(r[1560], c[1666], r[1668], c[1668]);
FA FA_1523(c[1442], r[1443], c[1560], r[1669], c[1669]);
FA FA_1524(r[1444], r[1445], c[1561], r[1670], c[1670]);
FA FA_1525(c[1445], r[1446], c[1563], r[1671], c[1671]);
FA FA_1526(c[1313], r[1314], c[1446], r[1672], c[1672]);
HA HA_146(r[1447], c[1564], r[1673], c[1673]);
FA FA_1527(c[1447], r[1448], c[1566], r[1674], c[1674]);
FA FA_1528(r[1316], r[1317], c[1448], r[1675], c[1675]);
HA HA_147(r[1449], c[1567], r[1676], c[1676]);
FA FA_1529(c[1449], r[1450], c[1569], r[1677], c[1677]);
FA FA_1530(r[1320], r[1321], r[1322], r[1678], c[1678]);
FA FA_1531(r[1323], r[1324], c[1451], r[1679], c[1679]);
HA HA_148(r[1452], r[1453], r[1680], c[1680]);
FA FA_1532(r[1327], c[1452], c[1453], r[1681], c[1681]);
FA FA_1533(r[1328], r[1329], c[1454], r[1682], c[1682]);
FA FA_1534(r[1331], c[1456], c[1457], r[1683], c[1683]);
FA FA_1535(c[1458], c[1459], c[1460], r[1684], c[1684]);
FA FA_1536(c[1462], r[1463], r[1464], r[1685], c[1685]);
FA FA_1537(c[1463], c[1464], c[1465], r[1686], c[1686]);
FA FA_1538(c[1467], r[1468], r[1469], r[1687], c[1687]);
FA FA_1539(c[1468], c[1469], c[1470], r[1688], c[1688]);
FA FA_1540(c[1472], r[1473], r[1474], r[1689], c[1689]);
FA FA_1541(c[1473], c[1474], c[1475], r[1690], c[1690]);
FA FA_1542(r[1476], r[1477], r[1478], r[1691], c[1691]);
FA FA_1543(c[1478], r[1479], r[1480], r[1692], c[1692]);
HA HA_149(r[1481], c[1590], r[1693], c[1693]);
FA FA_1544(c[1479], c[1480], c[1481], r[1694], c[1694]);
FA FA_1545(r[1482], r[1483], r[1484], r[1695], c[1695]);
FA FA_1546(c[1484], r[1485], r[1486], r[1696], c[1696]);
HA HA_150(r[1487], c[1595], r[1697], c[1697]);
FA FA_1547(r[1355], c[1485], c[1486], r[1698], c[1698]);
FA FA_1548(c[1487], r[1488], r[1489], r[1699], c[1699]);
HA HA_151(c[1597], c[1598], r[1700], c[1700]);
FA FA_1549(r[1358], c[1488], c[1489], r[1701], c[1701]);
FA FA_1550(r[1490], r[1491], r[1492], r[1702], c[1702]);
HA HA_152(c[1600], c[1601], r[1703], c[1703]);
FA FA_1551(r[1360], r[1361], c[1490], r[1704], c[1704]);
FA FA_1552(c[1491], c[1492], r[1493], r[1705], c[1705]);
FA FA_1553(r[1363], r[1364], c[1493], r[1706], c[1706]);
FA FA_1554(c[1494], r[1495], r[1496], r[1707], c[1707]);
HA HA_153(c[1605], c[1606], r[1708], c[1708]);
FA FA_1555(r[1366], r[1367], c[1495], r[1709], c[1709]);
FA FA_1556(c[1496], r[1497], r[1498], r[1710], c[1710]);
FA FA_1557(r[1369], r[1370], c[1497], r[1711], c[1711]);
FA FA_1558(c[1498], r[1499], r[1500], r[1712], c[1712]);
HA HA_154(c[1611], c[1612], r[1713], c[1713]);
FA FA_1559(c[1370], r[1371], r[1372], r[1714], c[1714]);
FA FA_1560(r[1373], c[1499], c[1500], r[1715], c[1715]);
HA HA_155(r[1501], r[1502], r[1716], c[1716]);
FA FA_1561(r[1375], r[1376], c[1501], r[1717], c[1717]);
FA FA_1562(c[1502], c[1503], r[1504], r[1718], c[1718]);
FA FA_1563(c[1376], r[1377], r[1378], r[1719], c[1719]);
FA FA_1564(r[1379], c[1504], c[1505], r[1720], c[1720]);
FA FA_1565(c[1379], r[1380], r[1381], r[1721], c[1721]);
FA FA_1566(r[1382], c[1506], c[1507], r[1722], c[1722]);
FA FA_1567(c[1382], r[1383], r[1384], r[1723], c[1723]);
FA FA_1568(r[1385], c[1509], c[1510], r[1724], c[1724]);
FA FA_1569(c[1385], r[1386], r[1387], r[1725], c[1725]);
FA FA_1570(r[1388], c[1512], c[1513], r[1726], c[1726]);
FA FA_1571(r[1389], r[1390], r[1391], r[1727], c[1727]);
FA FA_1572(r[1392], c[1515], c[1516], r[1728], c[1728]);
FA FA_1573(c[1392], r[1393], r[1394], r[1729], c[1729]);
FA FA_1574(r[1395], c[1518], c[1519], r[1730], c[1730]);
HA HA_156(c[1520], r[1521], r[1731], c[1731]);
FA FA_1575(c[1395], r[1396], r[1397], r[1732], c[1732]);
FA FA_1576(r[1398], c[1521], c[1522], r[1733], c[1733]);
FA FA_1577(r[1399], r[1400], r[1401], r[1734], c[1734]);
FA FA_1578(r[1402], c[1524], c[1525], r[1735], c[1735]);
HA HA_157(c[1526], r[1527], r[1736], c[1736]);
FA FA_1579(r[1403], r[1404], r[1405], r[1737], c[1737]);
FA FA_1580(r[1406], c[1527], c[1528], r[1738], c[1738]);
FA FA_1581(r[1407], r[1408], r[1409], r[1739], c[1739]);
FA FA_1582(r[1410], c[1530], c[1531], r[1740], c[1740]);
FA FA_1583(r[1411], r[1412], r[1413], r[1741], c[1741]);
FA FA_1584(r[1414], c[1533], c[1534], r[1742], c[1742]);
FA FA_1585(r[1415], r[1416], r[1417], r[1743], c[1743]);
FA FA_1586(r[1418], c[1536], c[1537], r[1744], c[1744]);
FA FA_1587(r[1421], r[1422], r[1423], r[1745], c[1745]);
FA FA_1588(c[1539], c[1540], c[1541], r[1746], c[1746]);
FA FA_1589(c[1423], r[1424], r[1425], r[1747], c[1747]);
FA FA_1590(r[1426], r[1427], c[1542], r[1748], c[1748]);
HA HA_158(c[1543], c[1544], r[1749], c[1749]);
HA HA_159(r[1661], r[1662], r[1750], c[1750]);
FA FA_1591(r[1557], c[1661], c[1662], r[1751], c[1751]);
HA HA_160(r[1663], c[1750], r[1752], c[1752]);
FA FA_1592(r[1664], r[1665], c[1751], r[1753], c[1753]);
FA FA_1593(r[1559], c[1664], c[1665], r[1754], c[1754]);
HA HA_161(r[1666], c[1753], r[1755], c[1755]);
FA FA_1594(r[1667], r[1668], c[1754], r[1756], c[1756]);
FA FA_1595(r[1561], r[1562], c[1667], r[1757], c[1757]);
FA FA_1596(c[1562], r[1563], c[1669], r[1758], c[1758]);
HA HA_162(r[1670], c[1757], r[1759], c[1759]);
FA FA_1597(r[1564], r[1565], c[1670], r[1760], c[1760]);
FA FA_1598(c[1565], r[1566], c[1671], r[1761], c[1761]);
FA FA_1599(r[1567], r[1568], c[1672], r[1762], c[1762]);
FA FA_1600(c[1568], r[1569], c[1674], r[1763], c[1763]);
FA FA_1601(r[1570], r[1571], c[1675], r[1764], c[1764]);
FA FA_1602(c[1450], r[1451], c[1570], r[1765], c[1765]);
HA HA_163(c[1571], r[1572], r[1766], c[1766]);
FA FA_1603(c[1572], r[1573], c[1678], r[1767], c[1767]);
FA FA_1604(r[1454], r[1455], c[1573], r[1768], c[1768]);
HA HA_164(r[1574], c[1679], r[1769], c[1769]);
FA FA_1605(c[1455], r[1456], r[1457], r[1770], c[1770]);
FA FA_1606(r[1458], r[1459], r[1460], r[1771], c[1771]);
HA HA_165(c[1575], r[1576], r[1772], c[1772]);
FA FA_1607(r[1461], r[1462], c[1576], r[1773], c[1773]);
FA FA_1608(r[1465], c[1577], c[1578], r[1774], c[1774]);
HA HA_166(r[1579], r[1580], r[1775], c[1775]);
FA FA_1609(r[1466], r[1467], c[1579], r[1776], c[1776]);
FA FA_1610(r[1470], c[1581], c[1582], r[1777], c[1777]);
HA HA_167(r[1583], r[1584], r[1778], c[1778]);
FA FA_1611(r[1471], r[1472], c[1583], r[1779], c[1779]);
FA FA_1612(r[1475], c[1585], c[1586], r[1780], c[1780]);
FA FA_1613(c[1587], c[1588], c[1589], r[1781], c[1781]);
FA FA_1614(c[1591], r[1592], r[1593], r[1782], c[1782]);
FA FA_1615(c[1592], c[1593], c[1594], r[1783], c[1783]);
FA FA_1616(c[1596], r[1597], r[1598], r[1784], c[1784]);
FA FA_1617(c[1599], r[1600], r[1601], r[1785], c[1785]);
FA FA_1618(c[1602], r[1603], r[1604], r[1786], c[1786]);
FA FA_1619(r[1494], c[1603], c[1604], r[1787], c[1787]);
FA FA_1620(r[1605], r[1606], r[1607], r[1788], c[1788]);
FA FA_1621(c[1607], r[1608], r[1609], r[1789], c[1789]);
HA HA_168(r[1610], c[1704], r[1790], c[1790]);
FA FA_1622(c[1608], c[1609], c[1610], r[1791], c[1791]);
FA FA_1623(r[1611], r[1612], r[1613], r[1792], c[1792]);
FA FA_1624(c[1613], r[1614], r[1615], r[1793], c[1793]);
HA HA_169(r[1616], c[1709], r[1794], c[1794]);
FA FA_1625(r[1503], c[1614], c[1615], r[1795], c[1795]);
FA FA_1626(c[1616], r[1617], r[1618], r[1796], c[1796]);
HA HA_170(c[1711], c[1712], r[1797], c[1797]);
FA FA_1627(r[1505], c[1617], c[1618], r[1798], c[1798]);
FA FA_1628(r[1619], r[1620], r[1621], r[1799], c[1799]);
HA HA_171(c[1714], c[1715], r[1800], c[1800]);
FA FA_1629(r[1506], r[1507], r[1508], r[1801], c[1801]);
FA FA_1630(c[1619], c[1620], c[1621], r[1802], c[1802]);
FA FA_1631(c[1508], r[1509], r[1510], r[1803], c[1803]);
FA FA_1632(r[1511], c[1622], c[1623], r[1804], c[1804]);
HA HA_172(r[1624], r[1625], r[1805], c[1805]);
FA FA_1633(c[1511], r[1512], r[1513], r[1806], c[1806]);
FA FA_1634(r[1514], c[1624], c[1625], r[1807], c[1807]);
FA FA_1635(c[1514], r[1515], r[1516], r[1808], c[1808]);
FA FA_1636(r[1517], c[1626], c[1627], r[1809], c[1809]);
HA HA_173(r[1628], r[1629], r[1810], c[1810]);
FA FA_1637(c[1517], r[1518], r[1519], r[1811], c[1811]);
FA FA_1638(r[1520], c[1628], c[1629], r[1812], c[1812]);
FA FA_1639(r[1522], r[1523], c[1630], r[1813], c[1813]);
FA FA_1640(c[1631], r[1632], r[1633], r[1814], c[1814]);
HA HA_174(r[1634], c[1727], r[1815], c[1815]);
FA FA_1641(c[1523], r[1524], r[1525], r[1816], c[1816]);
FA FA_1642(r[1526], c[1632], c[1633], r[1817], c[1817]);
FA FA_1643(r[1528], r[1529], c[1635], r[1818], c[1818]);
FA FA_1644(c[1636], c[1637], r[1638], r[1819], c[1819]);
HA HA_175(r[1639], c[1732], r[1820], c[1820]);
FA FA_1645(c[1529], r[1530], r[1531], r[1821], c[1821]);
FA FA_1646(r[1532], c[1638], c[1639], r[1822], c[1822]);
HA HA_176(r[1640], r[1641], r[1823], c[1823]);
FA FA_1647(c[1532], r[1533], r[1534], r[1824], c[1824]);
FA FA_1648(r[1535], c[1640], c[1641], r[1825], c[1825]);
HA HA_177(c[1642], r[1643], r[1826], c[1826]);
FA FA_1649(c[1535], r[1536], r[1537], r[1827], c[1827]);
FA FA_1650(r[1538], c[1643], c[1644], r[1828], c[1828]);
HA HA_178(c[1645], r[1646], r[1829], c[1829]);
FA FA_1651(c[1538], r[1539], r[1540], r[1830], c[1830]);
FA FA_1652(r[1541], c[1646], c[1647], r[1831], c[1831]);
HA HA_179(c[1648], r[1649], r[1832], c[1832]);
FA FA_1653(r[1542], r[1543], r[1544], r[1833], c[1833]);
FA FA_1654(r[1545], c[1649], c[1650], r[1834], c[1834]);
HA HA_180(c[1651], r[1652], r[1835], c[1835]);
FA FA_1655(c[1545], r[1546], r[1547], r[1836], c[1836]);
FA FA_1656(r[1548], c[1652], c[1653], r[1837], c[1837]);
HA HA_181(r[1751], r[1752], r[1838], c[1838]);
FA FA_1657(c[1752], r[1753], c[1838], r[1839], c[1839]);
FA FA_1658(r[1754], r[1755], c[1839], r[1840], c[1840]);
FA FA_1659(c[1755], r[1756], c[1840], r[1841], c[1841]);
FA FA_1660(c[1668], r[1669], c[1756], r[1842], c[1842]);
HA HA_182(r[1757], c[1841], r[1843], c[1843]);
FA FA_1661(r[1758], r[1759], c[1842], r[1844], c[1844]);
FA FA_1662(r[1671], c[1758], c[1759], r[1845], c[1845]);
HA HA_183(r[1760], c[1844], r[1846], c[1846]);
FA FA_1663(r[1672], r[1673], c[1760], r[1847], c[1847]);
FA FA_1664(c[1673], r[1674], c[1761], r[1848], c[1848]);
HA HA_184(r[1762], c[1847], r[1849], c[1849]);
FA FA_1665(r[1675], r[1676], c[1762], r[1850], c[1850]);
FA FA_1666(c[1676], r[1677], c[1763], r[1851], c[1851]);
HA HA_185(r[1764], c[1850], r[1852], c[1852]);
FA FA_1667(c[1677], r[1678], c[1764], r[1853], c[1853]);
FA FA_1668(r[1679], r[1680], c[1765], r[1854], c[1854]);
FA FA_1669(c[1680], r[1681], c[1767], r[1855], c[1855]);
FA FA_1670(c[1574], r[1575], c[1681], r[1856], c[1856]);
HA HA_186(r[1682], c[1768], r[1857], c[1857]);
FA FA_1671(c[1682], r[1683], c[1770], r[1858], c[1858]);
FA FA_1672(r[1577], r[1578], c[1683], r[1859], c[1859]);
HA HA_187(r[1684], c[1771], r[1860], c[1860]);
FA FA_1673(c[1684], r[1685], c[1773], r[1861], c[1861]);
FA FA_1674(c[1580], r[1581], r[1582], r[1862], c[1862]);
FA FA_1675(c[1686], r[1687], c[1776], r[1863], c[1863]);
FA FA_1676(c[1584], r[1585], r[1586], r[1864], c[1864]);
FA FA_1677(r[1587], r[1588], r[1589], r[1865], c[1865]);
HA HA_188(c[1688], r[1689], r[1866], c[1866]);
FA FA_1678(r[1590], r[1591], c[1689], r[1867], c[1867]);
FA FA_1679(r[1594], c[1690], c[1691], r[1868], c[1868]);
HA HA_189(r[1692], r[1693], r[1869], c[1869]);
FA FA_1680(r[1595], r[1596], c[1692], r[1870], c[1870]);
FA FA_1681(r[1599], c[1694], c[1695], r[1871], c[1871]);
HA HA_190(r[1696], r[1697], r[1872], c[1872]);
FA FA_1682(r[1602], c[1696], c[1697], r[1873], c[1873]);
FA FA_1683(c[1698], c[1699], c[1700], r[1874], c[1874]);
FA FA_1684(c[1701], c[1702], c[1703], r[1875], c[1875]);
FA FA_1685(c[1705], r[1706], r[1707], r[1876], c[1876]);
FA FA_1686(c[1706], c[1707], c[1708], r[1877], c[1877]);
FA FA_1687(c[1710], r[1711], r[1712], r[1878], c[1878]);
FA FA_1688(c[1713], r[1714], r[1715], r[1879], c[1879]);
FA FA_1689(c[1716], r[1717], r[1718], r[1880], c[1880]);
FA FA_1690(r[1622], r[1623], c[1717], r[1881], c[1881]);
FA FA_1691(c[1718], r[1719], r[1720], r[1882], c[1882]);
FA FA_1692(c[1719], c[1720], r[1721], r[1883], c[1883]);
HA HA_191(r[1722], c[1801], r[1884], c[1884]);
FA FA_1693(r[1626], r[1627], c[1721], r[1885], c[1885]);
FA FA_1694(c[1722], r[1723], r[1724], r[1886], c[1886]);
FA FA_1695(c[1723], c[1724], r[1725], r[1887], c[1887]);
HA HA_192(r[1726], c[1806], r[1888], c[1888]);
FA FA_1696(r[1630], r[1631], c[1725], r[1889], c[1889]);
FA FA_1697(c[1726], r[1727], r[1728], r[1890], c[1890]);
FA FA_1698(c[1728], r[1729], r[1730], r[1891], c[1891]);
HA HA_193(r[1731], c[1811], r[1892], c[1892]);
FA FA_1699(c[1634], r[1635], r[1636], r[1893], c[1893]);
FA FA_1700(r[1637], c[1729], c[1730], r[1894], c[1894]);
FA FA_1701(c[1733], r[1734], r[1735], r[1895], c[1895]);
HA HA_194(r[1736], c[1816], r[1896], c[1896]);
FA FA_1702(r[1642], c[1734], c[1735], r[1897], c[1897]);
FA FA_1703(c[1736], r[1737], r[1738], r[1898], c[1898]);
HA HA_195(c[1818], c[1819], r[1899], c[1899]);
FA FA_1704(r[1644], r[1645], c[1737], r[1900], c[1900]);
FA FA_1705(c[1738], r[1739], r[1740], r[1901], c[1901]);
FA FA_1706(r[1647], r[1648], c[1739], r[1902], c[1902]);
FA FA_1707(c[1740], r[1741], r[1742], r[1903], c[1903]);
HA HA_196(c[1824], c[1825], r[1904], c[1904]);
FA FA_1708(r[1650], r[1651], c[1741], r[1905], c[1905]);
FA FA_1709(c[1742], r[1743], r[1744], r[1906], c[1906]);
FA FA_1710(r[1653], r[1654], c[1743], r[1907], c[1907]);
FA FA_1711(c[1744], r[1745], r[1746], r[1908], c[1908]);
HA HA_197(c[1830], c[1831], r[1909], c[1909]);
FA FA_1712(c[1654], r[1655], r[1656], r[1910], c[1910]);
FA FA_1713(r[1657], c[1745], c[1746], r[1911], c[1911]);
HA HA_198(r[1747], r[1748], r[1912], c[1912]);
HA HA_199(r[1842], r[1843], r[1913], c[1913]);
FA FA_1714(c[1843], r[1844], c[1913], r[1914], c[1914]);
FA FA_1715(r[1845], r[1846], c[1914], r[1915], c[1915]);
FA FA_1716(r[1761], c[1845], c[1846], r[1916], c[1916]);
HA HA_200(r[1847], c[1915], r[1917], c[1917]);
FA FA_1717(r[1848], r[1849], c[1916], r[1918], c[1918]);
FA FA_1718(r[1763], c[1848], c[1849], r[1919], c[1919]);
HA HA_201(r[1850], c[1918], r[1920], c[1920]);
FA FA_1719(r[1851], r[1852], c[1919], r[1921], c[1921]);
FA FA_1720(r[1765], r[1766], c[1851], r[1922], c[1922]);
FA FA_1721(c[1766], r[1767], c[1853], r[1923], c[1923]);
HA HA_202(r[1854], c[1922], r[1924], c[1924]);
FA FA_1722(r[1768], r[1769], c[1854], r[1925], c[1925]);
FA FA_1723(c[1769], r[1770], c[1855], r[1926], c[1926]);
FA FA_1724(r[1771], r[1772], c[1856], r[1927], c[1927]);
FA FA_1725(c[1772], r[1773], c[1858], r[1928], c[1928]);
FA FA_1726(r[1774], r[1775], c[1859], r[1929], c[1929]);
FA FA_1727(c[1685], r[1686], c[1774], r[1930], c[1930]);
HA HA_203(c[1775], r[1776], r[1931], c[1931]);
FA FA_1728(r[1777], r[1778], c[1862], r[1932], c[1932]);
FA FA_1729(c[1687], r[1688], c[1777], r[1933], c[1933]);
HA HA_204(c[1778], r[1779], r[1934], c[1934]);
FA FA_1730(c[1779], r[1780], c[1864], r[1935], c[1935]);
FA FA_1731(r[1690], r[1691], c[1780], r[1936], c[1936]);
HA HA_205(r[1781], c[1865], r[1937], c[1937]);
FA FA_1732(c[1781], r[1782], c[1867], r[1938], c[1938]);
FA FA_1733(c[1693], r[1694], r[1695], r[1939], c[1939]);
FA FA_1734(c[1783], r[1784], c[1870], r[1940], c[1940]);
FA FA_1735(r[1698], r[1699], r[1700], r[1941], c[1941]);
FA FA_1736(r[1701], r[1702], r[1703], r[1942], c[1942]);
HA HA_206(c[1785], r[1786], r[1943], c[1943]);
FA FA_1737(r[1704], r[1705], c[1786], r[1944], c[1944]);
FA FA_1738(r[1708], c[1787], c[1788], r[1945], c[1945]);
HA HA_207(r[1789], r[1790], r[1946], c[1946]);
FA FA_1739(r[1709], r[1710], c[1789], r[1947], c[1947]);
FA FA_1740(r[1713], c[1791], c[1792], r[1948], c[1948]);
HA HA_208(r[1793], r[1794], r[1949], c[1949]);
FA FA_1741(r[1716], c[1793], c[1794], r[1950], c[1950]);
FA FA_1742(c[1795], c[1796], c[1797], r[1951], c[1951]);
FA FA_1743(c[1798], c[1799], c[1800], r[1952], c[1952]);
FA FA_1744(c[1802], r[1803], r[1804], r[1953], c[1953]);
FA FA_1745(c[1803], c[1804], c[1805], r[1954], c[1954]);
FA FA_1746(c[1807], r[1808], r[1809], r[1955], c[1955]);
FA FA_1747(c[1808], c[1809], c[1810], r[1956], c[1956]);
FA FA_1748(c[1812], r[1813], r[1814], r[1957], c[1957]);
FA FA_1749(c[1731], r[1732], r[1733], r[1958], c[1958]);
FA FA_1750(c[1813], c[1814], c[1815], r[1959], c[1959]);
FA FA_1751(c[1817], r[1818], r[1819], r[1960], c[1960]);
FA FA_1752(c[1820], r[1821], r[1822], r[1961], c[1961]);
FA FA_1753(c[1821], c[1822], c[1823], r[1962], c[1962]);
FA FA_1754(r[1824], r[1825], r[1826], r[1963], c[1963]);
FA FA_1755(c[1826], r[1827], r[1828], r[1964], c[1964]);
HA HA_209(r[1829], c[1900], r[1965], c[1965]);
FA FA_1756(c[1827], c[1828], c[1829], r[1966], c[1966]);
FA FA_1757(r[1830], r[1831], r[1832], r[1967], c[1967]);
FA FA_1758(c[1832], r[1833], r[1834], r[1968], c[1968]);
HA HA_210(r[1835], c[1905], r[1969], c[1969]);
FA FA_1759(r[1749], c[1833], c[1834], r[1970], c[1970]);
FA FA_1760(c[1835], r[1836], r[1837], r[1971], c[1971]);
HA HA_211(c[1907], c[1908], r[1972], c[1972]);
HA HA_212(r[1916], r[1917], r[1973], c[1973]);
FA FA_1761(c[1917], r[1918], c[1973], r[1974], c[1974]);
FA FA_1762(r[1919], r[1920], c[1974], r[1975], c[1975]);
FA FA_1763(c[1920], r[1921], c[1975], r[1976], c[1976]);
FA FA_1764(c[1852], r[1853], c[1921], r[1977], c[1977]);
HA HA_213(r[1922], c[1976], r[1978], c[1978]);
FA FA_1765(r[1923], r[1924], c[1977], r[1979], c[1979]);
FA FA_1766(r[1855], c[1923], c[1924], r[1980], c[1980]);
HA HA_214(r[1925], c[1979], r[1981], c[1981]);
FA FA_1767(r[1856], r[1857], c[1925], r[1982], c[1982]);
FA FA_1768(c[1857], r[1858], c[1926], r[1983], c[1983]);
HA HA_215(r[1927], c[1982], r[1984], c[1984]);
FA FA_1769(r[1859], r[1860], c[1927], r[1985], c[1985]);
FA FA_1770(c[1860], r[1861], c[1928], r[1986], c[1986]);
HA HA_216(r[1929], c[1985], r[1987], c[1987]);
FA FA_1771(c[1861], r[1862], c[1929], r[1988], c[1988]);
FA FA_1772(r[1863], c[1930], c[1931], r[1989], c[1989]);
HA HA_217(r[1932], c[1988], r[1990], c[1990]);
FA FA_1773(c[1863], r[1864], c[1932], r[1991], c[1991]);
FA FA_1774(r[1865], r[1866], c[1933], r[1992], c[1992]);
FA FA_1775(c[1866], r[1867], c[1935], r[1993], c[1993]);
FA FA_1776(r[1868], r[1869], c[1936], r[1994], c[1994]);
FA FA_1777(c[1782], r[1783], c[1868], r[1995], c[1995]);
HA HA_218(c[1869], r[1870], r[1996], c[1996]);
FA FA_1778(r[1871], r[1872], c[1939], r[1997], c[1997]);
FA FA_1779(c[1784], r[1785], c[1871], r[1998], c[1998]);
HA HA_219(c[1872], r[1873], r[1999], c[1999]);
FA FA_1780(c[1873], r[1874], c[1941], r[2000], c[2000]);
FA FA_1781(r[1787], r[1788], c[1874], r[2001], c[2001]);
HA HA_220(r[1875], c[1942], r[2002], c[2002]);
FA FA_1782(c[1875], r[1876], c[1944], r[2003], c[2003]);
FA FA_1783(c[1790], r[1791], r[1792], r[2004], c[2004]);
FA FA_1784(c[1877], r[1878], c[1947], r[2005], c[2005]);
FA FA_1785(r[1795], r[1796], r[1797], r[2006], c[2006]);
FA FA_1786(r[1798], r[1799], r[1800], r[2007], c[2007]);
HA HA_221(c[1879], r[1880], r[2008], c[2008]);
FA FA_1787(r[1801], r[1802], c[1880], r[2009], c[2009]);
FA FA_1788(r[1805], c[1881], c[1882], r[2010], c[2010]);
HA HA_222(r[1883], r[1884], r[2011], c[2011]);
FA FA_1789(r[1806], r[1807], c[1883], r[2012], c[2012]);
FA FA_1790(r[1810], c[1885], c[1886], r[2013], c[2013]);
HA HA_223(r[1887], r[1888], r[2014], c[2014]);
FA FA_1791(r[1811], r[1812], c[1887], r[2015], c[2015]);
FA FA_1792(r[1815], c[1889], c[1890], r[2016], c[2016]);
HA HA_224(r[1891], r[1892], r[2017], c[2017]);
FA FA_1793(r[1816], r[1817], c[1891], r[2018], c[2018]);
HA HA_225(c[1892], r[1893], r[2019], c[2019]);
FA FA_1794(r[1820], c[1893], c[1894], r[2020], c[2020]);
FA FA_1795(r[1823], c[1895], c[1896], r[2021], c[2021]);
FA FA_1796(c[1897], c[1898], c[1899], r[2022], c[2022]);
FA FA_1797(c[1901], r[1902], r[1903], r[2023], c[2023]);
FA FA_1798(c[1902], c[1903], c[1904], r[2024], c[2024]);
FA FA_1799(c[1906], r[1907], r[1908], r[2025], c[2025]);
FA FA_1800(c[1909], r[1910], r[1911], r[2026], c[2026]);
HA HA_226(r[1977], r[1978], r[2027], c[2027]);
FA FA_1801(c[1978], r[1979], c[2027], r[2028], c[2028]);
FA FA_1802(r[1980], r[1981], c[2028], r[2029], c[2029]);
FA FA_1803(r[1926], c[1980], c[1981], r[2030], c[2030]);
HA HA_227(r[1982], c[2029], r[2031], c[2031]);
FA FA_1804(r[1983], r[1984], c[2030], r[2032], c[2032]);
FA FA_1805(r[1928], c[1983], c[1984], r[2033], c[2033]);
HA HA_228(r[1985], c[2032], r[2034], c[2034]);
FA FA_1806(r[1986], r[1987], c[2033], r[2035], c[2035]);
FA FA_1807(r[1930], r[1931], c[1986], r[2036], c[2036]);
FA FA_1808(r[1989], r[1990], c[2036], r[2037], c[2037]);
FA FA_1809(r[1933], r[1934], c[1989], r[2038], c[2038]);
FA FA_1810(c[1934], r[1935], c[1991], r[2039], c[2039]);
HA HA_229(r[1992], c[2038], r[2040], c[2040]);
FA FA_1811(r[1936], r[1937], c[1992], r[2041], c[2041]);
FA FA_1812(c[1937], r[1938], c[1993], r[2042], c[2042]);
HA HA_230(r[1994], c[2041], r[2043], c[2043]);
FA FA_1813(c[1938], r[1939], c[1994], r[2044], c[2044]);
FA FA_1814(r[1940], c[1995], c[1996], r[2045], c[2045]);
HA HA_231(r[1997], c[2044], r[2046], c[2046]);
FA FA_1815(c[1940], r[1941], c[1997], r[2047], c[2047]);
FA FA_1816(r[1942], r[1943], c[1998], r[2048], c[2048]);
FA FA_1817(c[1943], r[1944], c[2000], r[2049], c[2049]);
FA FA_1818(r[1945], r[1946], c[2001], r[2050], c[2050]);
FA FA_1819(c[1876], r[1877], c[1945], r[2051], c[2051]);
HA HA_232(c[1946], r[1947], r[2052], c[2052]);
FA FA_1820(r[1948], r[1949], c[2004], r[2053], c[2053]);
FA FA_1821(c[1878], r[1879], c[1948], r[2054], c[2054]);
HA HA_233(c[1949], r[1950], r[2055], c[2055]);
FA FA_1822(c[1950], r[1951], c[2006], r[2056], c[2056]);
FA FA_1823(r[1881], r[1882], c[1951], r[2057], c[2057]);
HA HA_234(r[1952], c[2007], r[2058], c[2058]);
FA FA_1824(c[1952], r[1953], c[2009], r[2059], c[2059]);
FA FA_1825(c[1884], r[1885], r[1886], r[2060], c[2060]);
FA FA_1826(c[1954], r[1955], c[2012], r[2061], c[2061]);
FA FA_1827(c[1888], r[1889], r[1890], r[2062], c[2062]);
FA FA_1828(c[1956], r[1957], c[2015], r[2063], c[2063]);
FA FA_1829(r[1894], c[1957], r[1958], r[2064], c[2064]);
FA FA_1830(r[1895], r[1896], c[1958], r[2065], c[2065]);
FA FA_1831(r[1897], r[1898], r[1899], r[2066], c[2066]);
HA HA_235(c[1960], r[1961], r[2067], c[2067]);
FA FA_1832(r[1900], r[1901], c[1961], r[2068], c[2068]);
FA FA_1833(r[1904], c[1962], c[1963], r[2069], c[2069]);
HA HA_236(r[1964], r[1965], r[2070], c[2070]);
FA FA_1834(r[1905], r[1906], c[1964], r[2071], c[2071]);
FA FA_1835(r[1909], c[1966], c[1967], r[2072], c[2072]);
HA HA_237(r[1968], r[1969], r[2073], c[2073]);
FA FA_1836(r[1912], c[1968], c[1969], r[2074], c[2074]);
HA HA_238(r[2030], r[2031], r[2075], c[2075]);
FA FA_1837(c[2031], r[2032], c[2075], r[2076], c[2076]);
FA FA_1838(r[2033], r[2034], c[2076], r[2077], c[2077]);
FA FA_1839(c[2034], r[2035], c[2077], r[2078], c[2078]);
FA FA_1840(c[1987], r[1988], c[2035], r[2079], c[2079]);
HA HA_239(r[2036], c[2078], r[2080], c[2080]);
FA FA_1841(r[2037], c[2079], c[2080], r[2081], c[2081]);
FA FA_1842(c[1990], r[1991], c[2037], r[2082], c[2082]);
HA HA_240(r[2038], c[2081], r[2083], c[2083]);
FA FA_1843(r[2039], r[2040], c[2082], r[2084], c[2084]);
FA FA_1844(r[1993], c[2039], c[2040], r[2085], c[2085]);
HA HA_241(r[2041], c[2084], r[2086], c[2086]);
FA FA_1845(r[2042], r[2043], c[2085], r[2087], c[2087]);
FA FA_1846(r[1995], r[1996], c[2042], r[2088], c[2088]);
FA FA_1847(r[2045], r[2046], c[2088], r[2089], c[2089]);
FA FA_1848(r[1998], r[1999], c[2045], r[2090], c[2090]);
FA FA_1849(c[1999], r[2000], c[2047], r[2091], c[2091]);
HA HA_242(r[2048], c[2090], r[2092], c[2092]);
FA FA_1850(r[2001], r[2002], c[2048], r[2093], c[2093]);
FA FA_1851(c[2002], r[2003], c[2049], r[2094], c[2094]);
HA HA_243(r[2050], c[2093], r[2095], c[2095]);
FA FA_1852(c[2003], r[2004], c[2050], r[2096], c[2096]);
FA FA_1853(r[2005], c[2051], c[2052], r[2097], c[2097]);
HA HA_244(r[2053], c[2096], r[2098], c[2098]);
FA FA_1854(c[2005], r[2006], c[2053], r[2099], c[2099]);
FA FA_1855(r[2007], r[2008], c[2054], r[2100], c[2100]);
FA FA_1856(c[2008], r[2009], c[2056], r[2101], c[2101]);
FA FA_1857(r[2010], r[2011], c[2057], r[2102], c[2102]);
FA FA_1858(c[1953], r[1954], c[2010], r[2103], c[2103]);
HA HA_245(c[2011], r[2012], r[2104], c[2104]);
FA FA_1859(r[2013], r[2014], c[2060], r[2105], c[2105]);
FA FA_1860(c[1955], r[1956], c[2013], r[2106], c[2106]);
HA HA_246(c[2014], r[2015], r[2107], c[2107]);
FA FA_1861(r[2016], r[2017], c[2062], r[2108], c[2108]);
FA FA_1862(r[1959], c[2016], c[2017], r[2109], c[2109]);
HA HA_247(r[2018], r[2019], r[2110], c[2110]);
FA FA_1863(c[1959], r[1960], c[2018], r[2111], c[2111]);
FA FA_1864(c[2020], r[2021], c[2065], r[2112], c[2112]);
FA FA_1865(r[1962], r[1963], c[2021], r[2113], c[2113]);
HA HA_248(r[2022], c[2066], r[2114], c[2114]);
FA FA_1866(c[2022], r[2023], c[2068], r[2115], c[2115]);
FA FA_1867(c[1965], r[1966], r[1967], r[2116], c[2116]);
FA FA_1868(c[2024], r[2025], c[2071], r[2117], c[2117]);
FA FA_1869(r[1970], r[1971], r[1972], r[2118], c[2118]);
HA HA_249(r[2079], r[2080], r[2119], c[2119]);
HA HA_250(r[2081], c[2119], r[2120], c[2120]);
FA FA_1870(r[2082], r[2083], c[2120], r[2121], c[2121]);
FA FA_1871(c[2083], r[2084], c[2121], r[2122], c[2122]);
FA FA_1872(r[2085], r[2086], c[2122], r[2123], c[2123]);
FA FA_1873(c[2086], r[2087], c[2123], r[2124], c[2124]);
FA FA_1874(c[2043], r[2044], c[2087], r[2125], c[2125]);
HA HA_251(r[2088], c[2124], r[2126], c[2126]);
FA FA_1875(r[2089], c[2125], c[2126], r[2127], c[2127]);
FA FA_1876(c[2046], r[2047], c[2089], r[2128], c[2128]);
HA HA_252(r[2090], c[2127], r[2129], c[2129]);
FA FA_1877(r[2091], r[2092], c[2128], r[2130], c[2130]);
FA FA_1878(r[2049], c[2091], c[2092], r[2131], c[2131]);
HA HA_253(r[2093], c[2130], r[2132], c[2132]);
FA FA_1879(r[2094], r[2095], c[2131], r[2133], c[2133]);
FA FA_1880(r[2051], r[2052], c[2094], r[2134], c[2134]);
FA FA_1881(r[2097], r[2098], c[2134], r[2135], c[2135]);
FA FA_1882(r[2054], r[2055], c[2097], r[2136], c[2136]);
FA FA_1883(c[2055], r[2056], c[2099], r[2137], c[2137]);
HA HA_254(r[2100], c[2136], r[2138], c[2138]);
FA FA_1884(r[2057], r[2058], c[2100], r[2139], c[2139]);
FA FA_1885(c[2058], r[2059], c[2101], r[2140], c[2140]);
HA HA_255(r[2102], c[2139], r[2141], c[2141]);
FA FA_1886(c[2059], r[2060], c[2102], r[2142], c[2142]);
FA FA_1887(r[2061], c[2103], c[2104], r[2143], c[2143]);
HA HA_256(r[2105], c[2142], r[2144], c[2144]);
FA FA_1888(c[2061], r[2062], c[2105], r[2145], c[2145]);
FA FA_1889(r[2063], c[2106], c[2107], r[2146], c[2146]);
HA HA_257(r[2108], c[2145], r[2147], c[2147]);
FA FA_1890(c[2063], r[2064], c[2108], r[2148], c[2148]);
FA FA_1891(c[2019], r[2020], c[2064], r[2149], c[2149]);
HA HA_258(r[2065], c[2109], r[2150], c[2150]);
FA FA_1892(r[2066], r[2067], c[2111], r[2151], c[2151]);
FA FA_1893(c[2067], r[2068], c[2112], r[2152], c[2152]);
FA FA_1894(r[2069], r[2070], c[2113], r[2153], c[2153]);
FA FA_1895(c[2023], r[2024], c[2069], r[2154], c[2154]);
HA HA_259(c[2070], r[2071], r[2155], c[2155]);
FA FA_1896(r[2072], r[2073], c[2116], r[2156], c[2156]);
FA FA_1897(c[2025], r[2026], c[2072], r[2157], c[2157]);
HA HA_260(c[2073], r[2074], r[2158], c[2158]);
HA HA_261(r[2125], r[2126], r[2159], c[2159]);
HA HA_262(r[2127], c[2159], r[2160], c[2160]);
FA FA_1898(r[2128], r[2129], c[2160], r[2161], c[2161]);
FA FA_1899(c[2129], r[2130], c[2161], r[2162], c[2162]);
FA FA_1900(r[2131], r[2132], c[2162], r[2163], c[2163]);
FA FA_1901(c[2132], r[2133], c[2163], r[2164], c[2164]);
FA FA_1902(c[2095], r[2096], c[2133], r[2165], c[2165]);
HA HA_263(r[2134], c[2164], r[2166], c[2166]);
FA FA_1903(r[2135], c[2165], c[2166], r[2167], c[2167]);
FA FA_1904(c[2098], r[2099], c[2135], r[2168], c[2168]);
HA HA_264(r[2136], c[2167], r[2169], c[2169]);
FA FA_1905(r[2137], r[2138], c[2168], r[2170], c[2170]);
FA FA_1906(r[2101], c[2137], c[2138], r[2171], c[2171]);
HA HA_265(r[2139], c[2170], r[2172], c[2172]);
FA FA_1907(r[2140], r[2141], c[2171], r[2173], c[2173]);
FA FA_1908(r[2103], r[2104], c[2140], r[2174], c[2174]);
FA FA_1909(r[2143], r[2144], c[2174], r[2175], c[2175]);
FA FA_1910(r[2106], r[2107], c[2143], r[2176], c[2176]);
FA FA_1911(r[2146], r[2147], c[2176], r[2177], c[2177]);
FA FA_1912(r[2109], r[2110], c[2146], r[2178], c[2178]);
FA FA_1913(c[2110], r[2111], c[2148], r[2179], c[2179]);
FA FA_1914(r[2112], c[2149], c[2150], r[2180], c[2180]);
HA HA_266(r[2151], c[2179], r[2181], c[2181]);
FA FA_1915(r[2113], r[2114], c[2151], r[2182], c[2182]);
FA FA_1916(c[2114], r[2115], c[2152], r[2183], c[2183]);
HA HA_267(r[2153], c[2182], r[2184], c[2184]);
FA FA_1917(c[2115], r[2116], c[2153], r[2185], c[2185]);
FA FA_1918(r[2117], c[2154], c[2155], r[2186], c[2186]);
HA HA_268(r[2156], c[2185], r[2187], c[2187]);
FA FA_1919(c[2117], r[2118], c[2156], r[2188], c[2188]);
HA HA_269(r[2165], r[2166], r[2189], c[2189]);
HA HA_270(r[2167], c[2189], r[2190], c[2190]);
FA FA_1920(r[2168], r[2169], c[2190], r[2191], c[2191]);
FA FA_1921(c[2169], r[2170], c[2191], r[2192], c[2192]);
FA FA_1922(r[2171], r[2172], c[2192], r[2193], c[2193]);
FA FA_1923(c[2172], r[2173], c[2193], r[2194], c[2194]);
FA FA_1924(c[2141], r[2142], c[2173], r[2195], c[2195]);
HA HA_271(r[2174], c[2194], r[2196], c[2196]);
FA FA_1925(r[2175], c[2195], c[2196], r[2197], c[2197]);
FA FA_1926(c[2144], r[2145], c[2175], r[2198], c[2198]);
HA HA_272(r[2176], c[2197], r[2199], c[2199]);
FA FA_1927(r[2177], c[2198], c[2199], r[2200], c[2200]);
FA FA_1928(c[2147], r[2148], c[2177], r[2201], c[2201]);
HA HA_273(r[2178], c[2200], r[2202], c[2202]);
FA FA_1929(r[2149], r[2150], c[2178], r[2203], c[2203]);
FA FA_1930(r[2180], r[2181], c[2203], r[2204], c[2204]);
FA FA_1931(r[2152], c[2180], c[2181], r[2205], c[2205]);
HA HA_274(r[2182], c[2204], r[2206], c[2206]);
FA FA_1932(r[2183], r[2184], c[2205], r[2207], c[2207]);
FA FA_1933(r[2154], r[2155], c[2183], r[2208], c[2208]);
FA FA_1934(r[2186], r[2187], c[2208], r[2209], c[2209]);
FA FA_1935(r[2157], r[2158], c[2186], r[2210], c[2210]);
HA HA_275(r[2195], r[2196], r[2211], c[2211]);
HA HA_276(r[2197], c[2211], r[2212], c[2212]);
FA FA_1936(r[2198], r[2199], c[2212], r[2213], c[2213]);
HA HA_277(r[2200], c[2213], r[2214], c[2214]);
FA FA_1937(r[2201], r[2202], c[2214], r[2215], c[2215]);
FA FA_1938(r[2179], c[2201], c[2202], r[2216], c[2216]);
HA HA_278(r[2203], c[2215], r[2217], c[2217]);
FA FA_1939(r[2204], c[2216], c[2217], r[2218], c[2218]);
FA FA_1940(r[2205], r[2206], c[2218], r[2219], c[2219]);
FA FA_1941(c[2206], r[2207], c[2219], r[2220], c[2220]);
FA FA_1942(c[2184], r[2185], c[2207], r[2221], c[2221]);
HA HA_279(r[2208], c[2220], r[2222], c[2222]);
FA FA_1943(r[2209], c[2221], c[2222], r[2223], c[2223]);
FA FA_1944(c[2187], r[2188], c[2209], r[2224], c[2224]);
HA HA_280(r[2210], c[2223], r[2225], c[2225]);
HA HA_281(r[2216], r[2217], r[2226], c[2226]);
HA HA_282(r[2218], c[2226], r[2227], c[2227]);
HA HA_283(r[2219], c[2227], r[2228], c[2228]);
HA HA_284(r[2220], c[2228], r[2229], c[2229]);
FA FA_1945(r[2221], r[2222], c[2229], r[2230], c[2230]);
HA HA_285(r[2223], c[2230], r[2231], c[2231]);
FA FA_1946(r[2224], r[2225], c[2231], r[2232], c[2232]);

assign result[0] = p[0][0];
assign result[1] = r[0];
assign result[2] = r[296];
assign result[3] = r[297];
assign result[4] = r[773];
assign result[5] = r[774];
assign result[6] = r[967];
assign result[7] = r[1293];
assign result[8] = r[1294];
assign result[9] = r[1428];
assign result[10] = r[1549];
assign result[11] = r[1550];
assign result[12] = r[1658];
assign result[13] = r[1659];
assign result[14] = r[1660];
assign result[15] = r[1750];
assign result[16] = r[1838];
assign result[17] = r[1839];
assign result[18] = r[1840];
assign result[19] = r[1841];
assign result[20] = r[1913];
assign result[21] = r[1914];
assign result[22] = r[1915];
assign result[23] = r[1973];
assign result[24] = r[1974];
assign result[25] = r[1975];
assign result[26] = r[1976];
assign result[27] = r[2027];
assign result[28] = r[2028];
assign result[29] = r[2029];
assign result[30] = r[2075];
assign result[31] = r[2076];
assign result[32] = r[2077];
assign result[33] = r[2078];
assign result[34] = r[2119];
assign result[35] = r[2120];
assign result[36] = r[2121];
assign result[37] = r[2122];
assign result[38] = r[2123];
assign result[39] = r[2124];
assign result[40] = r[2159];
assign result[41] = r[2160];
assign result[42] = r[2161];
assign result[43] = r[2162];
assign result[44] = r[2163];
assign result[45] = r[2164];
assign result[46] = r[2189];
assign result[47] = r[2190];
assign result[48] = r[2191];
assign result[49] = r[2192];
assign result[50] = r[2193];
assign result[51] = r[2194];
assign result[52] = r[2211];
assign result[53] = r[2212];
assign result[54] = r[2213];
assign result[55] = r[2214];
assign result[56] = r[2215];
assign result[57] = r[2226];
assign result[58] = r[2227];
assign result[59] = r[2228];
assign result[60] = r[2229];
assign result[61] = r[2230];
assign result[62] = r[2231];
assign result[63] = r[2232];

endmodule

module registerNbits #(
    parameter N = 8
) (
    clk,
    reset,
    en,
    inp,
    out
);
  input clk, reset, en;
  output reg [N-1:0] out;
  input [N-1:0] inp;
  always @(posedge clk) begin
    if (reset) out <= 'b0;
    else if (en) out <= inp;

  end
endmodule


module signed_wallace (
    input i_clk,
    input i_rst,
    input i_en,
    input [31:0] i_inputA,
    input [31:0] i_inputB,
    output [63:0] o_result
);

  wire [31:0] A_reg;
  wire [31:0] B_reg;
  wire [63:0] out_reg;


  registerNbits #(32) regA (
      i_clk,
      i_rst,
      i_en,
      i_inputA,
      A_reg
  );
  registerNbits #(32) regB (
      i_clk,
      i_rst,
      i_en,
      i_inputB,
      B_reg
  );
  signed_wallace_tree_multipler unt (
      A_reg,
      B_reg,
      out_reg
  );
  registerNbits #(64) outReg (
      i_clk,
      i_rst,
      i_en,
      out_reg,
      o_result[63:0]
  );


endmodule