/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Dec 20 14:16:31 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2098498826 */

module n_case(A, B, S, outA, outB, enable);
   input [31:0]A;
   input [31:0]B;
   output [31:0]S;
   output [2:0]outA;
   output [2:0]outB;
   output enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_4;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;

   AND2_X1 i_0_0 (.A1(outB[0]), .A2(outA[0]), .ZN(enable));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_0), .ZN(S[22]));
   OAI22_X1 i_0_2 (.A1(outB[1]), .A2(outB[0]), .B1(outA[1]), .B2(outA[0]), 
      .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(S[30]));
   OAI22_X1 i_0_4 (.A1(n_0_21), .A2(outA[2]), .B1(n_0_16), .B2(outB[2]), 
      .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .ZN(S[31]));
   XNOR2_X1 i_0_6 (.A(B[31]), .B(A[31]), .ZN(n_0_2));
   AOI22_X1 i_0_7 (.A1(outA[2]), .A2(n_0_5), .B1(n_0_7), .B2(outB[2]), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_21), .A2(n_0_17), .ZN(n_0_5));
   AOI21_X1 i_0_9 (.A(outA[2]), .B1(n_0_28), .B2(n_0_17), .ZN(outA[0]));
   AOI21_X1 i_0_10 (.A(n_0_28), .B1(n_0_17), .B2(outA[2]), .ZN(outA[1]));
   NOR2_X1 i_0_11 (.A1(n_0_20), .A2(n_0_19), .ZN(outA[2]));
   NAND4_X1 i_0_12 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_0_19));
   NAND4_X1 i_0_13 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(outB[2]), .B1(n_0_31), .B2(n_0_8), .ZN(outB[0]));
   NAND2_X1 i_0_15 (.A1(n_0_31), .A2(n_0_8), .ZN(n_0_21));
   AOI21_X1 i_0_16 (.A(n_0_31), .B1(n_0_8), .B2(outB[2]), .ZN(outB[1]));
   AND2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_32), .ZN(n_0_31));
   NOR4_X1 i_0_18 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_32));
   NOR4_X1 i_0_19 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_33));
   NOR2_X1 i_0_20 (.A1(n_0_6), .A2(n_0_4), .ZN(outB[2]));
   NAND4_X1 i_0_21 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_4));
   NAND4_X1 i_0_22 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_0_6));
   NAND2_X1 i_0_23 (.A1(n_0_16), .A2(n_0_8), .ZN(n_0_7));
   AND3_X1 i_0_24 (.A1(n_0_10), .A2(n_0_9), .A3(n_0_11), .ZN(n_0_8));
   NOR4_X1 i_0_25 (.A1(B[19]), .A2(B[18]), .A3(B[16]), .A4(B[12]), .ZN(n_0_9));
   NOR4_X1 i_0_26 (.A1(B[17]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n_0_10));
   NOR4_X1 i_0_27 (.A1(B[10]), .A2(B[9]), .A3(B[8]), .A4(n_0_12), .ZN(n_0_11));
   NAND3_X1 i_0_28 (.A1(n_0_14), .A2(n_0_13), .A3(n_0_15), .ZN(n_0_12));
   NOR4_X1 i_0_29 (.A1(B[5]), .A2(B[3]), .A3(B[2]), .A4(B[1]), .ZN(n_0_13));
   NOR4_X1 i_0_30 (.A1(B[22]), .A2(B[21]), .A3(B[20]), .A4(B[0]), .ZN(n_0_14));
   NOR4_X1 i_0_31 (.A1(B[11]), .A2(B[7]), .A3(B[6]), .A4(B[4]), .ZN(n_0_15));
   NAND2_X1 i_0_32 (.A1(n_0_28), .A2(n_0_17), .ZN(n_0_16));
   AND3_X1 i_0_33 (.A1(n_0_22), .A2(n_0_18), .A3(n_0_23), .ZN(n_0_17));
   NOR4_X1 i_0_34 (.A1(A[19]), .A2(A[18]), .A3(A[16]), .A4(A[12]), .ZN(n_0_18));
   NOR4_X1 i_0_35 (.A1(A[17]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n_0_22));
   NOR4_X1 i_0_36 (.A1(A[10]), .A2(A[9]), .A3(A[8]), .A4(n_0_24), .ZN(n_0_23));
   NAND3_X1 i_0_37 (.A1(n_0_26), .A2(n_0_25), .A3(n_0_27), .ZN(n_0_24));
   NOR4_X1 i_0_38 (.A1(A[5]), .A2(A[3]), .A3(A[2]), .A4(A[1]), .ZN(n_0_25));
   NOR4_X1 i_0_39 (.A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[0]), .ZN(n_0_26));
   NOR4_X1 i_0_40 (.A1(A[11]), .A2(A[7]), .A3(A[6]), .A4(A[4]), .ZN(n_0_27));
   AND2_X1 i_0_41 (.A1(n_0_30), .A2(n_0_29), .ZN(n_0_28));
   NOR4_X1 i_0_42 (.A1(A[25]), .A2(A[24]), .A3(A[30]), .A4(A[27]), .ZN(n_0_29));
   NOR4_X1 i_0_43 (.A1(A[26]), .A2(A[23]), .A3(A[29]), .A4(A[28]), .ZN(n_0_30));
endmodule

module zero_counter(M, Zcount);
   input [23:0]M;
   output [4:0]Zcount;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_0), .B2(Zcount[4]), .ZN(Zcount[0]));
   OAI21_X1 i_0_1 (.A(n_0_33), .B1(M[6]), .B2(n_0_1), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(M[5]), .A2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(M[4]), .A2(n_0_3), .ZN(n_0_2));
   NOR2_X1 i_0_4 (.A1(M[3]), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(M[2]), .B1(n_0_32), .B2(M[0]), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(n_0_6), .B1(n_0_9), .B2(n_0_27), .ZN(n_0_5));
   AOI211_X1 i_0_7 (.A(M[15]), .B(n_0_27), .C1(n_0_7), .C2(n_0_36), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_35), .B1(M[12]), .B2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(M[11]), .B1(n_0_34), .B2(M[9]), .ZN(n_0_8));
   AOI221_X1 i_0_10 (.A(M[23]), .B1(n_0_39), .B2(M[21]), .C1(n_0_30), .C2(n_0_10), 
      .ZN(n_0_9));
   OAI21_X1 i_0_11 (.A(n_0_38), .B1(n_0_37), .B2(M[18]), .ZN(n_0_10));
   AOI21_X1 i_0_12 (.A(n_0_14), .B1(n_0_11), .B2(Zcount[4]), .ZN(Zcount[1]));
   OR3_X1 i_0_13 (.A1(M[7]), .A2(M[6]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(M[5]), .A2(M[4]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(M[3]), .A2(M[2]), .A3(n_0_23), .ZN(n_0_13));
   AOI22_X1 i_0_16 (.A1(n_0_26), .A2(n_0_17), .B1(n_0_15), .B2(n_0_27), .ZN(
      n_0_14));
   NOR3_X1 i_0_17 (.A1(M[23]), .A2(M[22]), .A3(n_0_16), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(M[21]), .A2(M[20]), .A3(n_0_29), .ZN(n_0_16));
   OAI21_X1 i_0_19 (.A(n_0_25), .B1(M[10]), .B2(M[11]), .ZN(n_0_17));
   OAI21_X1 i_0_20 (.A(n_0_18), .B1(n_0_19), .B2(Zcount[4]), .ZN(Zcount[2]));
   NAND3_X1 i_0_21 (.A1(Zcount[4]), .A2(n_0_22), .A3(n_0_21), .ZN(n_0_18));
   AOI22_X1 i_0_22 (.A1(n_0_26), .A2(n_0_25), .B1(n_0_30), .B2(n_0_27), .ZN(
      n_0_19));
   OAI22_X1 i_0_23 (.A1(n_0_22), .A2(n_0_20), .B1(n_0_27), .B2(Zcount[4]), 
      .ZN(Zcount[3]));
   NAND2_X1 i_0_24 (.A1(Zcount[4]), .A2(n_0_21), .ZN(n_0_20));
   NOR4_X1 i_0_25 (.A1(M[7]), .A2(M[6]), .A3(M[5]), .A4(M[4]), .ZN(n_0_21));
   NAND2_X1 i_0_26 (.A1(n_0_24), .A2(n_0_23), .ZN(n_0_22));
   NOR2_X1 i_0_27 (.A1(M[1]), .A2(M[0]), .ZN(n_0_23));
   NOR2_X1 i_0_28 (.A1(M[3]), .A2(M[2]), .ZN(n_0_24));
   AND3_X1 i_0_29 (.A1(n_0_31), .A2(n_0_26), .A3(n_0_25), .ZN(Zcount[4]));
   NOR2_X1 i_0_30 (.A1(M[13]), .A2(M[12]), .ZN(n_0_25));
   NOR3_X1 i_0_31 (.A1(n_0_27), .A2(M[14]), .A3(M[15]), .ZN(n_0_26));
   NAND3_X1 i_0_32 (.A1(n_0_30), .A2(n_0_29), .A3(n_0_28), .ZN(n_0_27));
   NOR2_X1 i_0_33 (.A1(M[17]), .A2(M[16]), .ZN(n_0_28));
   NOR2_X1 i_0_34 (.A1(M[19]), .A2(M[18]), .ZN(n_0_29));
   NOR4_X1 i_0_35 (.A1(M[23]), .A2(M[22]), .A3(M[21]), .A4(M[20]), .ZN(n_0_30));
   NOR4_X1 i_0_36 (.A1(M[11]), .A2(M[10]), .A3(M[9]), .A4(M[8]), .ZN(n_0_31));
   INV_X1 i_0_37 (.A(M[1]), .ZN(n_0_32));
   INV_X1 i_0_38 (.A(M[7]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(M[10]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(M[13]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(M[14]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(M[17]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(M[19]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(M[22]), .ZN(n_0_39));
endmodule

module datapath__0_29(Nb, Na, mult_res);
   input [23:0]Nb;
   input [23:0]Na;
   output [47:0]mult_res;

   HA_X1 i_0 (.A(n_1538), .B(n_1694), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(n_1514), .B(n_1537), .CI(n_1560), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(n_1581), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(n_1559), .B(n_1580), .CI(n_5), .CO(n_8), .S(n_6));
   FA_X1 i_4 (.A(n_1466), .B(n_1489), .CI(n_1512), .CO(n_13), .S(n_9));
   FA_X1 i_5 (.A(n_1535), .B(n_1558), .CI(n_1579), .CO(n_15), .S(n_10));
   FA_X1 i_6 (.A(n_1442), .B(n_1465), .CI(n_1488), .CO(n_21), .S(n_12));
   FA_X1 i_7 (.A(n_1511), .B(n_1534), .CI(n_1557), .CO(n_23), .S(n_14));
   FA_X1 i_8 (.A(n_1578), .B(n_15), .CI(n_13), .CO(n_25), .S(n_20));
   FA_X1 i_9 (.A(n_1418), .B(n_1441), .CI(n_1464), .CO(n_31), .S(n_22));
   FA_X1 i_10 (.A(n_1487), .B(n_1510), .CI(n_1533), .CO(n_33), .S(n_24));
   FA_X1 i_11 (.A(n_1556), .B(n_1577), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_12 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_32), .S(n_30));
   FA_X1 i_13 (.A(n_1394), .B(n_1417), .CI(n_1440), .CO(n_43), .S(n_42));
   FA_X1 i_14 (.A(n_1463), .B(n_1486), .CI(n_1509), .CO(n_45), .S(n_44));
   FA_X1 i_15 (.A(n_1532), .B(n_1555), .CI(n_1576), .CO(n_47), .S(n_46));
   FA_X1 i_16 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_36));
   FA_X1 i_17 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_48), .S(n_37));
   FA_X1 i_18 (.A(n_1370), .B(n_1393), .CI(n_1416), .CO(n_57), .S(n_56));
   FA_X1 i_19 (.A(n_1439), .B(n_1462), .CI(n_1485), .CO(n_59), .S(n_58));
   FA_X1 i_20 (.A(n_1508), .B(n_1531), .CI(n_1554), .CO(n_61), .S(n_60));
   FA_X1 i_21 (.A(n_1575), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_22 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_50));
   FA_X1 i_23 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_64), .S(n_51));
   FA_X1 i_24 (.A(n_1346), .B(n_1369), .CI(n_1392), .CO(n_73), .S(n_72));
   FA_X1 i_25 (.A(n_1415), .B(n_1438), .CI(n_1461), .CO(n_75), .S(n_74));
   FA_X1 i_26 (.A(n_1484), .B(n_1507), .CI(n_1530), .CO(n_77), .S(n_76));
   FA_X1 i_27 (.A(n_1553), .B(n_1574), .CI(n_61), .CO(n_66), .S(n_78));
   FA_X1 i_28 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_67), .S(n_80));
   FA_X1 i_29 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_81), .S(n_79));
   FA_X1 i_30 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_83), .S(n_82));
   FA_X1 i_45 (.A(n_1322), .B(n_1345), .CI(n_1368), .CO(n_85), .S(n_84));
   FA_X1 i_46 (.A(n_1391), .B(n_1414), .CI(n_1437), .CO(n_91), .S(n_90));
   FA_X1 i_47 (.A(n_1460), .B(n_1483), .CI(n_1506), .CO(n_95), .S(n_92));
   FA_X1 i_48 (.A(n_1529), .B(n_1552), .CI(n_1573), .CO(n_97), .S(n_93));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_96), .S(n_94));
   FA_X1 i_31 (.A(n_1298), .B(n_1321), .CI(n_1344), .CO(n_99), .S(n_98));
   FA_X1 i_56 (.A(n_1367), .B(n_1390), .CI(n_1413), .CO(n_111), .S(n_110));
   FA_X1 i_57 (.A(n_1436), .B(n_1459), .CI(n_1482), .CO(n_113), .S(n_112));
   FA_X1 i_32 (.A(n_1505), .B(n_1528), .CI(n_1551), .CO(n_117), .S(n_114));
   FA_X1 i_33 (.A(n_1572), .B(n_97), .CI(n_95), .CO(n_116), .S(n_115));
   FA_X1 i_34 (.A(n_1274), .B(n_1297), .CI(n_1320), .CO(n_133), .S(n_118));
   FA_X1 i_35 (.A(n_1343), .B(n_1366), .CI(n_1389), .CO(n_135), .S(n_119));
   FA_X1 i_36 (.A(n_1412), .B(n_1435), .CI(n_1458), .CO(n_137), .S(n_132));
   FA_X1 i_37 (.A(n_1481), .B(n_1504), .CI(n_1527), .CO(n_139), .S(n_134));
   FA_X1 i_38 (.A(n_1550), .B(n_1571), .CI(n_117), .CO(n_141), .S(n_136));
   FA_X1 i_39 (.A(n_1250), .B(n_1273), .CI(n_1296), .CO(n_140), .S(n_138));
   FA_X1 i_40 (.A(n_1319), .B(n_1342), .CI(n_1365), .CO(n_156), .S(n_143));
   FA_X1 i_41 (.A(n_1388), .B(n_1411), .CI(n_1434), .CO(n_158), .S(n_157));
   FA_X1 i_42 (.A(n_1457), .B(n_1480), .CI(n_1503), .CO(n_160), .S(n_159));
   FA_X1 i_43 (.A(n_1526), .B(n_1549), .CI(n_1570), .CO(n_162), .S(n_161));
   FA_X1 i_44 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_164), .S(n_163));
   FA_X1 i_50 (.A(n_133), .B(n_879), .CI(n_141), .CO(n_166), .S(n_165));
   FA_X1 i_51 (.A(n_1032), .B(n_1055), .CI(n_1078), .CO(n_167), .S(n_550));
   FA_X1 i_52 (.A(n_1101), .B(n_1124), .CI(n_1147), .CO(n_553), .S(n_552));
   FA_X1 i_53 (.A(n_1170), .B(n_1193), .CI(n_1216), .CO(n_555), .S(n_554));
   FA_X1 i_54 (.A(n_1239), .B(n_1262), .CI(n_1285), .CO(n_557), .S(n_556));
   FA_X1 i_55 (.A(n_1308), .B(n_1331), .CI(n_1354), .CO(n_559), .S(n_558));
   FA_X1 i_58 (.A(n_1377), .B(n_1400), .CI(n_1423), .CO(n_561), .S(n_560));
   FA_X1 i_59 (.A(n_1446), .B(n_1469), .CI(n_1492), .CO(n_563), .S(n_562));
   FA_X1 i_60 (.A(n_1515), .B(n_732), .CI(n_733), .CO(n_168), .S(n_564));
   FA_X1 i_61 (.A(n_698), .B(n_699), .CI(n_704), .CO(n_461), .S(n_169));
   FA_X1 i_62 (.A(n_694), .B(n_696), .CI(n_686), .CO(n_505), .S(n_504));
   FA_X1 i_63 (.A(n_688), .B(n_726), .CI(n_562), .CO(n_509), .S(n_507));
   FA_X1 i_64 (.A(n_560), .B(n_558), .CI(n_556), .CO(n_513), .S(n_511));
   FA_X1 i_65 (.A(n_554), .B(n_552), .CI(n_550), .CO(n_517), .S(n_515));
   FA_X1 i_66 (.A(n_564), .B(n_705), .CI(n_738), .CO(n_521), .S(n_519));
   FA_X1 i_67 (.A(n_1031), .B(n_1054), .CI(n_1077), .CO(n_525), .S(n_523));
   FA_X1 i_68 (.A(n_1100), .B(n_1123), .CI(n_1146), .CO(n_529), .S(n_527));
   FA_X1 i_69 (.A(n_1169), .B(n_1192), .CI(n_1215), .CO(n_533), .S(n_531));
   FA_X1 i_70 (.A(n_1238), .B(n_1261), .CI(n_1284), .CO(n_537), .S(n_535));
   FA_X1 i_71 (.A(n_1307), .B(n_1330), .CI(n_1353), .CO(n_541), .S(n_539));
   FA_X1 i_72 (.A(n_1376), .B(n_1399), .CI(n_1422), .CO(n_545), .S(n_543));
   FA_X1 i_73 (.A(n_1445), .B(n_1468), .CI(n_1491), .CO(n_548), .S(n_547));
   FA_X1 i_74 (.A(n_563), .B(n_561), .CI(n_559), .CO(n_551), .S(n_549));
   FA_X1 i_75 (.A(n_557), .B(n_555), .CI(n_553), .CO(n_566), .S(n_565));
   FA_X1 i_76 (.A(n_1726), .B(n_1728), .CI(n_1729), .CO(n_693), .S(n_567));
   FA_X1 i_77 (.A(n_1730), .B(n_1751), .CI(n_1736), .CO(n_569), .S(n_568));
   FA_X1 i_78 (.A(n_1737), .B(n_1752), .CI(n_1738), .CO(n_571), .S(n_570));
   FA_X1 i_79 (.A(n_693), .B(n_1731), .CI(n_1727), .CO(n_573), .S(n_572));
   FA_X1 i_80 (.A(n_1021), .B(n_1044), .CI(n_1067), .CO(n_903), .S(n_902));
   FA_X1 i_81 (.A(n_1090), .B(n_1113), .CI(n_1136), .CO(n_905), .S(n_904));
   FA_X1 i_82 (.A(n_1159), .B(n_1182), .CI(n_1205), .CO(n_907), .S(n_906));
   FA_X1 i_83 (.A(n_1228), .B(n_1251), .CI(n_1755), .CO(n_909), .S(n_908));
   FA_X1 i_84 (.A(n_1758), .B(n_1759), .CI(n_1760), .CO(n_911), .S(n_910));
   FA_X1 i_85 (.A(n_1762), .B(n_908), .CI(n_906), .CO(n_913), .S(n_912));
   FA_X1 i_86 (.A(n_904), .B(n_902), .CI(n_910), .CO(n_915), .S(n_914));
   FA_X1 i_87 (.A(n_1761), .B(n_1756), .CI(n_1769), .CO(n_917), .S(n_916));
   FA_X1 i_88 (.A(n_914), .B(n_912), .CI(n_1757), .CO(n_919), .S(n_918));
   FA_X1 i_89 (.A(n_916), .B(n_1770), .CI(n_918), .CO(n_921), .S(n_920));
   FA_X1 i_90 (.A(n_1020), .B(n_1043), .CI(n_1066), .CO(n_923), .S(n_922));
   FA_X1 i_91 (.A(n_1089), .B(n_1112), .CI(n_1135), .CO(n_925), .S(n_924));
   FA_X1 i_92 (.A(n_1158), .B(n_1181), .CI(n_1204), .CO(n_927), .S(n_926));
   FA_X1 i_93 (.A(n_1227), .B(n_907), .CI(n_905), .CO(n_929), .S(n_928));
   FA_X1 i_94 (.A(n_903), .B(n_911), .CI(n_909), .CO(n_931), .S(n_930));
   FA_X1 i_95 (.A(n_926), .B(n_924), .CI(n_922), .CO(n_933), .S(n_932));
   FA_X1 i_96 (.A(n_928), .B(n_913), .CI(n_930), .CO(n_935), .S(n_934));
   FA_X1 i_97 (.A(n_915), .B(n_932), .CI(n_917), .CO(n_937), .S(n_936));
   FA_X1 i_98 (.A(n_934), .B(n_919), .CI(n_936), .CO(n_939), .S(n_938));
   FA_X1 i_99 (.A(n_1019), .B(n_1042), .CI(n_1065), .CO(n_941), .S(n_940));
   FA_X1 i_100 (.A(n_1088), .B(n_1111), .CI(n_1134), .CO(n_943), .S(n_942));
   FA_X1 i_101 (.A(n_1157), .B(n_1180), .CI(n_1203), .CO(n_945), .S(n_944));
   FA_X1 i_102 (.A(n_927), .B(n_925), .CI(n_923), .CO(n_947), .S(n_946));
   FA_X1 i_103 (.A(n_929), .B(n_944), .CI(n_942), .CO(n_949), .S(n_948));
   FA_X1 i_104 (.A(n_940), .B(n_931), .CI(n_946), .CO(n_951), .S(n_950));
   FA_X1 i_105 (.A(n_933), .B(n_948), .CI(n_950), .CO(n_953), .S(n_952));
   FA_X1 i_106 (.A(n_935), .B(n_937), .CI(n_952), .CO(n_955), .S(n_954));
   FA_X1 i_107 (.A(n_1018), .B(n_1041), .CI(n_1064), .CO(n_957), .S(n_956));
   FA_X1 i_108 (.A(n_1087), .B(n_1110), .CI(n_1133), .CO(n_959), .S(n_958));
   FA_X1 i_109 (.A(n_1156), .B(n_1179), .CI(n_945), .CO(n_961), .S(n_960));
   FA_X1 i_110 (.A(n_943), .B(n_941), .CI(n_947), .CO(n_963), .S(n_962));
   FA_X1 i_111 (.A(n_960), .B(n_958), .CI(n_956), .CO(n_965), .S(n_964));
   FA_X1 i_112 (.A(n_962), .B(n_949), .CI(n_951), .CO(n_967), .S(n_966));
   FA_X1 i_113 (.A(n_964), .B(n_966), .CI(n_953), .CO(n_969), .S(n_968));
   FA_X1 i_114 (.A(n_1017), .B(n_1040), .CI(n_1063), .CO(n_971), .S(n_970));
   FA_X1 i_115 (.A(n_1086), .B(n_1109), .CI(n_1132), .CO(n_973), .S(n_972));
   FA_X1 i_116 (.A(n_1155), .B(n_959), .CI(n_957), .CO(n_975), .S(n_974));
   FA_X1 i_117 (.A(n_961), .B(n_972), .CI(n_970), .CO(n_977), .S(n_976));
   FA_X1 i_118 (.A(n_963), .B(n_974), .CI(n_965), .CO(n_979), .S(n_978));
   FA_X1 i_119 (.A(n_976), .B(n_967), .CI(n_978), .CO(n_981), .S(n_980));
   FA_X1 i_120 (.A(n_1016), .B(n_1039), .CI(n_1062), .CO(n_983), .S(n_982));
   FA_X1 i_121 (.A(n_1085), .B(n_1108), .CI(n_1131), .CO(n_985), .S(n_984));
   FA_X1 i_122 (.A(n_973), .B(n_971), .CI(n_975), .CO(n_987), .S(n_986));
   FA_X1 i_123 (.A(n_984), .B(n_982), .CI(n_986), .CO(n_989), .S(n_988));
   FA_X1 i_124 (.A(n_977), .B(n_979), .CI(n_988), .CO(n_991), .S(n_990));
   FA_X1 i_125 (.A(n_1015), .B(n_1038), .CI(n_1061), .CO(n_993), .S(n_992));
   FA_X1 i_126 (.A(n_1084), .B(n_1107), .CI(n_985), .CO(n_995), .S(n_994));
   FA_X1 i_127 (.A(n_983), .B(n_994), .CI(n_992), .CO(n_997), .S(n_996));
   FA_X1 i_128 (.A(n_987), .B(n_989), .CI(n_996), .CO(n_999), .S(n_998));
   FA_X1 i_129 (.A(n_1014), .B(n_1037), .CI(n_1060), .CO(n_1001), .S(n_1000));
   FA_X1 i_130 (.A(n_1083), .B(n_993), .CI(n_995), .CO(n_1003), .S(n_1002));
   FA_X1 i_131 (.A(n_1000), .B(n_1002), .CI(n_997), .CO(n_1005), .S(n_1004));
   FA_X1 i_132 (.A(n_1013), .B(n_1036), .CI(n_1059), .CO(n_1007), .S(n_1006));
   FA_X1 i_133 (.A(n_1001), .B(n_1006), .CI(n_1003), .CO(n_1009), .S(n_1008));
   FA_X1 i_134 (.A(n_1012), .B(n_1035), .CI(n_1007), .CO(n_1011), .S(n_1010));
   NOR2_X1 i_135 (.A1(n_1725), .A2(n_1699), .ZN(n_1012));
   NOR2_X1 i_136 (.A1(n_1725), .A2(n_1698), .ZN(n_1013));
   NOR2_X1 i_137 (.A1(n_1725), .A2(n_1697), .ZN(n_1014));
   NOR2_X1 i_138 (.A1(n_1725), .A2(n_1696), .ZN(n_1015));
   NOR2_X1 i_139 (.A1(n_1725), .A2(n_1691), .ZN(n_1016));
   NOR2_X1 i_140 (.A1(n_1725), .A2(n_1690), .ZN(n_1017));
   NOR2_X1 i_141 (.A1(n_1725), .A2(n_1689), .ZN(n_1018));
   NOR2_X1 i_142 (.A1(n_1725), .A2(n_1688), .ZN(n_1019));
   NOR2_X1 i_143 (.A1(n_1725), .A2(n_1687), .ZN(n_1020));
   NOR2_X1 i_144 (.A1(n_1725), .A2(n_1686), .ZN(n_1021));
   NOR2_X1 i_145 (.A1(n_1725), .A2(n_1674), .ZN(n_574));
   NOR2_X1 i_146 (.A1(n_1725), .A2(n_1673), .ZN(n_1031));
   NOR2_X1 i_147 (.A1(n_1725), .A2(n_1670), .ZN(n_1032));
   NOR2_X1 i_148 (.A1(n_1724), .A2(n_1700), .ZN(n_1035));
   NOR2_X1 i_149 (.A1(n_1724), .A2(n_1699), .ZN(n_1036));
   NOR2_X1 i_150 (.A1(n_1724), .A2(n_1698), .ZN(n_1037));
   NOR2_X1 i_151 (.A1(n_1724), .A2(n_1697), .ZN(n_1038));
   NOR2_X1 i_152 (.A1(n_1724), .A2(n_1696), .ZN(n_1039));
   NOR2_X1 i_153 (.A1(n_1724), .A2(n_1691), .ZN(n_1040));
   NOR2_X1 i_154 (.A1(n_1724), .A2(n_1690), .ZN(n_1041));
   NOR2_X1 i_155 (.A1(n_1724), .A2(n_1689), .ZN(n_1042));
   NOR2_X1 i_156 (.A1(n_1724), .A2(n_1688), .ZN(n_1043));
   NOR2_X1 i_157 (.A1(n_1724), .A2(n_1687), .ZN(n_1044));
   NOR2_X1 i_158 (.A1(n_1724), .A2(n_1676), .ZN(n_575));
   NOR2_X1 i_159 (.A1(n_1724), .A2(n_1674), .ZN(n_1054));
   NOR2_X1 i_160 (.A1(n_1724), .A2(n_1673), .ZN(n_1055));
   NOR2_X1 i_161 (.A1(n_1723), .A2(n_1700), .ZN(n_1059));
   NOR2_X1 i_162 (.A1(n_1723), .A2(n_1699), .ZN(n_1060));
   NOR2_X1 i_163 (.A1(n_1723), .A2(n_1698), .ZN(n_1061));
   NOR2_X1 i_164 (.A1(n_1723), .A2(n_1697), .ZN(n_1062));
   NOR2_X1 i_165 (.A1(n_1723), .A2(n_1696), .ZN(n_1063));
   NOR2_X1 i_166 (.A1(n_1723), .A2(n_1691), .ZN(n_1064));
   NOR2_X1 i_167 (.A1(n_1723), .A2(n_1690), .ZN(n_1065));
   NOR2_X1 i_168 (.A1(n_1723), .A2(n_1689), .ZN(n_1066));
   NOR2_X1 i_169 (.A1(n_1723), .A2(n_1688), .ZN(n_1067));
   NOR2_X1 i_170 (.A1(n_1723), .A2(n_1678), .ZN(n_578));
   NOR2_X1 i_171 (.A1(n_1723), .A2(n_1676), .ZN(n_1077));
   NOR2_X1 i_172 (.A1(n_1723), .A2(n_1674), .ZN(n_1078));
   NOR2_X1 i_173 (.A1(n_1722), .A2(n_1700), .ZN(n_1083));
   NOR2_X1 i_174 (.A1(n_1722), .A2(n_1699), .ZN(n_1084));
   NOR2_X1 i_175 (.A1(n_1722), .A2(n_1698), .ZN(n_1085));
   NOR2_X1 i_176 (.A1(n_1722), .A2(n_1697), .ZN(n_1086));
   NOR2_X1 i_177 (.A1(n_1722), .A2(n_1696), .ZN(n_1087));
   NOR2_X1 i_178 (.A1(n_1722), .A2(n_1691), .ZN(n_1088));
   NOR2_X1 i_179 (.A1(n_1722), .A2(n_1690), .ZN(n_1089));
   NOR2_X1 i_180 (.A1(n_1722), .A2(n_1689), .ZN(n_1090));
   NOR2_X1 i_181 (.A1(n_1722), .A2(n_1679), .ZN(n_579));
   NOR2_X1 i_182 (.A1(n_1722), .A2(n_1678), .ZN(n_1100));
   NOR2_X1 i_183 (.A1(n_1722), .A2(n_1676), .ZN(n_1101));
   NOR2_X1 i_184 (.A1(n_1721), .A2(n_1700), .ZN(n_1107));
   NOR2_X1 i_185 (.A1(n_1721), .A2(n_1699), .ZN(n_1108));
   NOR2_X1 i_186 (.A1(n_1721), .A2(n_1698), .ZN(n_1109));
   NOR2_X1 i_187 (.A1(n_1721), .A2(n_1697), .ZN(n_1110));
   NOR2_X1 i_188 (.A1(n_1721), .A2(n_1696), .ZN(n_1111));
   NOR2_X1 i_189 (.A1(n_1721), .A2(n_1691), .ZN(n_1112));
   NOR2_X1 i_190 (.A1(n_1721), .A2(n_1690), .ZN(n_1113));
   NOR2_X1 i_191 (.A1(n_1721), .A2(n_1681), .ZN(n_590));
   NOR2_X1 i_192 (.A1(n_1721), .A2(n_1679), .ZN(n_1123));
   NOR2_X1 i_193 (.A1(n_1721), .A2(n_1678), .ZN(n_1124));
   NOR2_X1 i_194 (.A1(n_1720), .A2(n_1700), .ZN(n_1131));
   NOR2_X1 i_195 (.A1(n_1720), .A2(n_1699), .ZN(n_1132));
   NOR2_X1 i_196 (.A1(n_1720), .A2(n_1698), .ZN(n_1133));
   NOR2_X1 i_197 (.A1(n_1720), .A2(n_1697), .ZN(n_1134));
   NOR2_X1 i_198 (.A1(n_1720), .A2(n_1696), .ZN(n_1135));
   NOR2_X1 i_199 (.A1(n_1720), .A2(n_1691), .ZN(n_1136));
   NOR2_X1 i_200 (.A1(n_1720), .A2(n_1682), .ZN(n_591));
   NOR2_X1 i_201 (.A1(n_1720), .A2(n_1681), .ZN(n_1146));
   NOR2_X1 i_202 (.A1(n_1720), .A2(n_1679), .ZN(n_1147));
   NOR2_X1 i_203 (.A1(n_1719), .A2(n_1700), .ZN(n_1155));
   NOR2_X1 i_204 (.A1(n_1719), .A2(n_1699), .ZN(n_1156));
   NOR2_X1 i_205 (.A1(n_1719), .A2(n_1698), .ZN(n_1157));
   NOR2_X1 i_206 (.A1(n_1719), .A2(n_1697), .ZN(n_1158));
   NOR2_X1 i_207 (.A1(n_1719), .A2(n_1696), .ZN(n_1159));
   NOR2_X1 i_208 (.A1(n_1719), .A2(n_1683), .ZN(n_592));
   NOR2_X1 i_209 (.A1(n_1719), .A2(n_1682), .ZN(n_1169));
   NOR2_X1 i_210 (.A1(n_1719), .A2(n_1681), .ZN(n_1170));
   NOR2_X1 i_211 (.A1(n_1718), .A2(n_1700), .ZN(n_1179));
   NOR2_X1 i_212 (.A1(n_1718), .A2(n_1699), .ZN(n_1180));
   NOR2_X1 i_213 (.A1(n_1718), .A2(n_1698), .ZN(n_1181));
   NOR2_X1 i_214 (.A1(n_1718), .A2(n_1697), .ZN(n_1182));
   NOR2_X1 i_215 (.A1(n_1718), .A2(n_1684), .ZN(n_593));
   NOR2_X1 i_216 (.A1(n_1718), .A2(n_1683), .ZN(n_1192));
   NOR2_X1 i_217 (.A1(n_1718), .A2(n_1682), .ZN(n_1193));
   NOR2_X1 i_218 (.A1(n_1716), .A2(n_1700), .ZN(n_1203));
   NOR2_X1 i_219 (.A1(n_1716), .A2(n_1699), .ZN(n_1204));
   NOR2_X1 i_220 (.A1(n_1716), .A2(n_1698), .ZN(n_1205));
   NOR2_X1 i_221 (.A1(n_1716), .A2(n_1685), .ZN(n_594));
   NOR2_X1 i_222 (.A1(n_1716), .A2(n_1684), .ZN(n_1215));
   NOR2_X1 i_223 (.A1(n_1716), .A2(n_1683), .ZN(n_1216));
   NOR2_X1 i_224 (.A1(n_1716), .A2(n_1615), .ZN(n_595));
   NOR2_X1 i_225 (.A1(n_1715), .A2(n_1700), .ZN(n_1227));
   NOR2_X1 i_226 (.A1(n_1715), .A2(n_1699), .ZN(n_1228));
   NOR2_X1 i_227 (.A1(n_1715), .A2(n_1686), .ZN(n_596));
   NOR2_X1 i_228 (.A1(n_1715), .A2(n_1685), .ZN(n_1238));
   NOR2_X1 i_229 (.A1(n_1715), .A2(n_1684), .ZN(n_1239));
   NOR2_X1 i_230 (.A1(n_1715), .A2(n_1669), .ZN(n_597));
   NOR2_X1 i_744 (.A1(n_1715), .A2(n_1615), .ZN(n_1250));
   NOR2_X1 i_231 (.A1(n_1714), .A2(n_1700), .ZN(n_1251));
   NOR2_X1 i_232 (.A1(n_1714), .A2(n_1687), .ZN(n_598));
   NOR2_X1 i_233 (.A1(n_1714), .A2(n_1686), .ZN(n_1261));
   NOR2_X1 i_234 (.A1(n_1714), .A2(n_1685), .ZN(n_1262));
   NOR2_X1 i_235 (.A1(n_1714), .A2(n_1670), .ZN(n_599));
   NOR2_X1 i_767 (.A1(n_1714), .A2(n_1669), .ZN(n_1273));
   NOR2_X1 i_236 (.A1(n_1714), .A2(n_1615), .ZN(n_1274));
   NOR2_X1 i_237 (.A1(n_1713), .A2(n_1688), .ZN(n_600));
   NOR2_X1 i_238 (.A1(n_1713), .A2(n_1687), .ZN(n_1284));
   NOR2_X1 i_239 (.A1(n_1713), .A2(n_1686), .ZN(n_1285));
   NOR2_X1 i_790 (.A1(n_1713), .A2(n_1670), .ZN(n_1296));
   NOR2_X1 i_240 (.A1(n_1713), .A2(n_1669), .ZN(n_1297));
   NOR2_X1 i_792 (.A1(n_1713), .A2(n_1615), .ZN(n_1298));
   NOR2_X1 i_241 (.A1(n_1712), .A2(n_1689), .ZN(n_601));
   NOR2_X1 i_242 (.A1(n_1712), .A2(n_1688), .ZN(n_1307));
   NOR2_X1 i_243 (.A1(n_1712), .A2(n_1687), .ZN(n_1308));
   NOR2_X1 i_813 (.A1(n_1712), .A2(n_1673), .ZN(n_1319));
   NOR2_X1 i_244 (.A1(n_1712), .A2(n_1670), .ZN(n_1320));
   NOR2_X1 i_815 (.A1(n_1712), .A2(n_1669), .ZN(n_1321));
   NOR2_X1 i_816 (.A1(n_1712), .A2(n_1615), .ZN(n_1322));
   NOR2_X1 i_245 (.A1(n_1711), .A2(n_1690), .ZN(n_602));
   NOR2_X1 i_246 (.A1(n_1711), .A2(n_1689), .ZN(n_1330));
   NOR2_X1 i_247 (.A1(n_1711), .A2(n_1688), .ZN(n_1331));
   NOR2_X1 i_836 (.A1(n_1711), .A2(n_1674), .ZN(n_1342));
   NOR2_X1 i_248 (.A1(n_1711), .A2(n_1673), .ZN(n_1343));
   NOR2_X1 i_838 (.A1(n_1711), .A2(n_1670), .ZN(n_1344));
   NOR2_X1 i_839 (.A1(n_1711), .A2(n_1669), .ZN(n_1345));
   NOR2_X1 i_249 (.A1(n_1711), .A2(n_1615), .ZN(n_1346));
   NOR2_X1 i_250 (.A1(n_1710), .A2(n_1691), .ZN(n_603));
   NOR2_X1 i_251 (.A1(n_1710), .A2(n_1690), .ZN(n_1353));
   NOR2_X1 i_252 (.A1(n_1710), .A2(n_1689), .ZN(n_1354));
   NOR2_X1 i_859 (.A1(n_1710), .A2(n_1676), .ZN(n_1365));
   NOR2_X1 i_253 (.A1(n_1710), .A2(n_1674), .ZN(n_1366));
   NOR2_X1 i_861 (.A1(n_1710), .A2(n_1673), .ZN(n_1367));
   NOR2_X1 i_862 (.A1(n_1710), .A2(n_1670), .ZN(n_1368));
   NOR2_X1 i_254 (.A1(n_1710), .A2(n_1669), .ZN(n_1369));
   NOR2_X1 i_255 (.A1(n_1710), .A2(n_1615), .ZN(n_1370));
   NOR2_X1 i_256 (.A1(n_1709), .A2(n_1696), .ZN(n_604));
   NOR2_X1 i_257 (.A1(n_1709), .A2(n_1691), .ZN(n_1376));
   NOR2_X1 i_258 (.A1(n_1709), .A2(n_1690), .ZN(n_1377));
   NOR2_X1 i_882 (.A1(n_1709), .A2(n_1678), .ZN(n_1388));
   NOR2_X1 i_259 (.A1(n_1709), .A2(n_1676), .ZN(n_1389));
   NOR2_X1 i_884 (.A1(n_1709), .A2(n_1674), .ZN(n_1390));
   NOR2_X1 i_885 (.A1(n_1709), .A2(n_1673), .ZN(n_1391));
   NOR2_X1 i_260 (.A1(n_1709), .A2(n_1670), .ZN(n_1392));
   NOR2_X1 i_261 (.A1(n_1709), .A2(n_1669), .ZN(n_1393));
   NOR2_X1 i_262 (.A1(n_1709), .A2(n_1615), .ZN(n_1394));
   NOR2_X1 i_263 (.A1(n_1708), .A2(n_1697), .ZN(n_605));
   NOR2_X1 i_264 (.A1(n_1708), .A2(n_1696), .ZN(n_1399));
   NOR2_X1 i_265 (.A1(n_1708), .A2(n_1691), .ZN(n_1400));
   NOR2_X1 i_905 (.A1(n_1708), .A2(n_1679), .ZN(n_1411));
   NOR2_X1 i_266 (.A1(n_1708), .A2(n_1678), .ZN(n_1412));
   NOR2_X1 i_907 (.A1(n_1708), .A2(n_1676), .ZN(n_1413));
   NOR2_X1 i_908 (.A1(n_1708), .A2(n_1674), .ZN(n_1414));
   NOR2_X1 i_267 (.A1(n_1708), .A2(n_1673), .ZN(n_1415));
   NOR2_X1 i_268 (.A1(n_1708), .A2(n_1670), .ZN(n_1416));
   NOR2_X1 i_269 (.A1(n_1708), .A2(n_1669), .ZN(n_1417));
   NOR2_X1 i_270 (.A1(n_1708), .A2(n_1615), .ZN(n_1418));
   NOR2_X1 i_271 (.A1(n_1707), .A2(n_1698), .ZN(n_606));
   NOR2_X1 i_272 (.A1(n_1707), .A2(n_1697), .ZN(n_1422));
   NOR2_X1 i_273 (.A1(n_1707), .A2(n_1696), .ZN(n_1423));
   NOR2_X1 i_928 (.A1(n_1707), .A2(n_1681), .ZN(n_1434));
   NOR2_X1 i_274 (.A1(n_1707), .A2(n_1679), .ZN(n_1435));
   NOR2_X1 i_930 (.A1(n_1707), .A2(n_1678), .ZN(n_1436));
   NOR2_X1 i_931 (.A1(n_1707), .A2(n_1676), .ZN(n_1437));
   NOR2_X1 i_275 (.A1(n_1707), .A2(n_1674), .ZN(n_1438));
   NOR2_X1 i_276 (.A1(n_1707), .A2(n_1673), .ZN(n_1439));
   NOR2_X1 i_277 (.A1(n_1707), .A2(n_1670), .ZN(n_1440));
   NOR2_X1 i_278 (.A1(n_1707), .A2(n_1669), .ZN(n_1441));
   NOR2_X1 i_279 (.A1(n_1707), .A2(n_1615), .ZN(n_1442));
   NOR2_X1 i_280 (.A1(n_1706), .A2(n_1699), .ZN(n_607));
   NOR2_X1 i_281 (.A1(n_1706), .A2(n_1698), .ZN(n_1445));
   NOR2_X1 i_282 (.A1(n_1706), .A2(n_1697), .ZN(n_1446));
   NOR2_X1 i_951 (.A1(n_1706), .A2(n_1682), .ZN(n_1457));
   NOR2_X1 i_283 (.A1(n_1706), .A2(n_1681), .ZN(n_1458));
   NOR2_X1 i_953 (.A1(n_1706), .A2(n_1679), .ZN(n_1459));
   NOR2_X1 i_954 (.A1(n_1706), .A2(n_1678), .ZN(n_1460));
   NOR2_X1 i_284 (.A1(n_1706), .A2(n_1676), .ZN(n_1461));
   NOR2_X1 i_285 (.A1(n_1706), .A2(n_1674), .ZN(n_1462));
   NOR2_X1 i_286 (.A1(n_1706), .A2(n_1673), .ZN(n_1463));
   NOR2_X1 i_287 (.A1(n_1706), .A2(n_1670), .ZN(n_1464));
   NOR2_X1 i_288 (.A1(n_1706), .A2(n_1669), .ZN(n_1465));
   NOR2_X1 i_289 (.A1(n_1706), .A2(n_1615), .ZN(n_1466));
   NOR2_X1 i_290 (.A1(n_1705), .A2(n_1700), .ZN(n_608));
   NOR2_X1 i_291 (.A1(n_1705), .A2(n_1699), .ZN(n_1468));
   NOR2_X1 i_292 (.A1(n_1705), .A2(n_1698), .ZN(n_1469));
   NOR2_X1 i_974 (.A1(n_1705), .A2(n_1683), .ZN(n_1480));
   NOR2_X1 i_293 (.A1(n_1705), .A2(n_1682), .ZN(n_1481));
   NOR2_X1 i_976 (.A1(n_1705), .A2(n_1681), .ZN(n_1482));
   NOR2_X1 i_977 (.A1(n_1705), .A2(n_1679), .ZN(n_1483));
   NOR2_X1 i_294 (.A1(n_1705), .A2(n_1678), .ZN(n_1484));
   NOR2_X1 i_295 (.A1(n_1705), .A2(n_1676), .ZN(n_1485));
   NOR2_X1 i_296 (.A1(n_1705), .A2(n_1674), .ZN(n_1486));
   NOR2_X1 i_297 (.A1(n_1705), .A2(n_1673), .ZN(n_1487));
   NOR2_X1 i_298 (.A1(n_1705), .A2(n_1670), .ZN(n_1488));
   NOR2_X1 i_299 (.A1(n_1705), .A2(n_1669), .ZN(n_1489));
   NOR2_X1 i_300 (.A1(n_1705), .A2(n_1615), .ZN(n_609));
   NOR2_X1 i_301 (.A1(n_1704), .A2(n_1700), .ZN(n_1491));
   NOR2_X1 i_302 (.A1(n_1704), .A2(n_1699), .ZN(n_1492));
   NOR2_X1 i_997 (.A1(n_1704), .A2(n_1684), .ZN(n_1503));
   NOR2_X1 i_303 (.A1(n_1704), .A2(n_1683), .ZN(n_1504));
   NOR2_X1 i_304 (.A1(n_1704), .A2(n_1682), .ZN(n_1505));
   NOR2_X1 i_1000 (.A1(n_1704), .A2(n_1681), .ZN(n_1506));
   NOR2_X1 i_305 (.A1(n_1704), .A2(n_1679), .ZN(n_1507));
   NOR2_X1 i_306 (.A1(n_1704), .A2(n_1678), .ZN(n_1508));
   NOR2_X1 i_307 (.A1(n_1704), .A2(n_1676), .ZN(n_1509));
   NOR2_X1 i_308 (.A1(n_1704), .A2(n_1674), .ZN(n_1510));
   NOR2_X1 i_309 (.A1(n_1704), .A2(n_1673), .ZN(n_1511));
   NOR2_X1 i_310 (.A1(n_1704), .A2(n_1670), .ZN(n_1512));
   NOR2_X1 i_311 (.A1(n_1704), .A2(n_1669), .ZN(n_630));
   NOR2_X1 i_312 (.A1(n_1704), .A2(n_1615), .ZN(n_1514));
   NOR2_X1 i_313 (.A1(n_1703), .A2(n_1700), .ZN(n_1515));
   NOR2_X1 i_1020 (.A1(n_1703), .A2(n_1685), .ZN(n_1526));
   NOR2_X1 i_314 (.A1(n_1703), .A2(n_1684), .ZN(n_1527));
   NOR2_X1 i_315 (.A1(n_1703), .A2(n_1683), .ZN(n_1528));
   NOR2_X1 i_1023 (.A1(n_1703), .A2(n_1682), .ZN(n_1529));
   NOR2_X1 i_316 (.A1(n_1703), .A2(n_1681), .ZN(n_1530));
   NOR2_X1 i_317 (.A1(n_1703), .A2(n_1679), .ZN(n_1531));
   NOR2_X1 i_318 (.A1(n_1703), .A2(n_1678), .ZN(n_1532));
   NOR2_X1 i_319 (.A1(n_1703), .A2(n_1676), .ZN(n_1533));
   NOR2_X1 i_320 (.A1(n_1703), .A2(n_1674), .ZN(n_1534));
   NOR2_X1 i_321 (.A1(n_1703), .A2(n_1673), .ZN(n_1535));
   NOR2_X1 i_322 (.A1(n_1703), .A2(n_1670), .ZN(n_631));
   NOR2_X1 i_323 (.A1(n_1703), .A2(n_1669), .ZN(n_1537));
   NOR2_X1 i_324 (.A1(n_1703), .A2(n_1615), .ZN(n_1538));
   NOR2_X1 i_1043 (.A1(n_1702), .A2(n_1686), .ZN(n_1549));
   NOR2_X1 i_325 (.A1(n_1702), .A2(n_1685), .ZN(n_1550));
   NOR2_X1 i_326 (.A1(n_1702), .A2(n_1684), .ZN(n_1551));
   NOR2_X1 i_1046 (.A1(n_1702), .A2(n_1683), .ZN(n_1552));
   NOR2_X1 i_327 (.A1(n_1702), .A2(n_1682), .ZN(n_1553));
   NOR2_X1 i_328 (.A1(n_1702), .A2(n_1681), .ZN(n_1554));
   NOR2_X1 i_329 (.A1(n_1702), .A2(n_1679), .ZN(n_1555));
   NOR2_X1 i_330 (.A1(n_1702), .A2(n_1678), .ZN(n_1556));
   NOR2_X1 i_331 (.A1(n_1702), .A2(n_1676), .ZN(n_1557));
   NOR2_X1 i_332 (.A1(n_1702), .A2(n_1674), .ZN(n_1558));
   NOR2_X1 i_1053 (.A1(n_1702), .A2(n_1673), .ZN(n_1559));
   NOR2_X1 i_333 (.A1(n_1702), .A2(n_1670), .ZN(n_1560));
   NOR2_X1 i_334 (.A1(n_1701), .A2(n_1688), .ZN(n_657));
   NOR2_X1 i_1064 (.A1(n_1701), .A2(n_1687), .ZN(n_1570));
   NOR2_X1 i_335 (.A1(n_1701), .A2(n_1686), .ZN(n_1571));
   NOR2_X1 i_1066 (.A1(n_1701), .A2(n_1685), .ZN(n_1572));
   NOR2_X1 i_1067 (.A1(n_1701), .A2(n_1684), .ZN(n_1573));
   NOR2_X1 i_336 (.A1(n_1701), .A2(n_1683), .ZN(n_1574));
   NOR2_X1 i_337 (.A1(n_1701), .A2(n_1682), .ZN(n_1575));
   NOR2_X1 i_338 (.A1(n_1701), .A2(n_1681), .ZN(n_1576));
   NOR2_X1 i_339 (.A1(n_1701), .A2(n_1679), .ZN(n_1577));
   NOR2_X1 i_340 (.A1(n_1701), .A2(n_1678), .ZN(n_1578));
   NOR2_X1 i_341 (.A1(n_1701), .A2(n_1676), .ZN(n_1579));
   NOR2_X1 i_1074 (.A1(n_1701), .A2(n_1674), .ZN(n_1580));
   NOR2_X1 i_342 (.A1(n_1701), .A2(n_1673), .ZN(n_1581));
   XOR2_X1 i_343 (.A(n_889), .B(n_1582), .Z(mult_res[23]));
   NOR2_X1 i_344 (.A1(n_1805), .A2(n_1583), .ZN(n_1582));
   XOR2_X1 i_345 (.A(n_1605), .B(n_1593), .Z(mult_res[25]));
   XOR2_X1 i_346 (.A(n_1592), .B(n_1589), .Z(mult_res[26]));
   XOR2_X1 i_347 (.A(n_1590), .B(n_1587), .Z(mult_res[27]));
   NOR2_X1 i_348 (.A1(n_668), .A2(n_1794), .ZN(n_1587));
   XNOR2_X1 i_349 (.A(n_1594), .B(n_1588), .ZN(mult_res[28]));
   OAI21_X1 i_350 (.A(n_1818), .B1(n_1794), .B2(n_1590), .ZN(n_1588));
   NOR2_X1 i_351 (.A1(n_669), .A2(n_1717), .ZN(n_1589));
   INV_X1 i_352 (.A(n_1591), .ZN(n_1590));
   OAI21_X1 i_353 (.A(n_1817), .B1(n_1717), .B2(n_1592), .ZN(n_1591));
   AOI21_X1 i_354 (.A(n_1802), .B1(n_1796), .B2(n_1605), .ZN(n_1592));
   OAI21_X1 i_355 (.A(n_1796), .B1(n_855), .B2(n_1747), .ZN(n_1593));
   AOI21_X1 i_356 (.A(n_670), .B1(n_1754), .B2(n_1744), .ZN(n_1594));
   XNOR2_X1 i_357 (.A(n_1604), .B(n_1603), .ZN(mult_res[29]));
   INV_X1 i_358 (.A(n_1595), .ZN(mult_res[30]));
   AOI21_X1 i_359 (.A(n_1599), .B1(n_1601), .B2(n_1600), .ZN(n_1595));
   XOR2_X1 i_360 (.A(n_1597), .B(n_1596), .Z(mult_res[31]));
   OAI21_X1 i_361 (.A(n_1811), .B1(n_1807), .B2(n_1601), .ZN(n_1596));
   OAI21_X1 i_362 (.A(n_1806), .B1(n_1743), .B2(n_1741), .ZN(n_1597));
   XNOR2_X1 i_363 (.A(n_1609), .B(n_1598), .ZN(mult_res[32]));
   OAI21_X1 i_364 (.A(n_1806), .B1(n_1810), .B2(n_1599), .ZN(n_1598));
   NOR2_X1 i_365 (.A1(n_1601), .A2(n_1600), .ZN(n_1599));
   OR2_X1 i_366 (.A1(n_1812), .A2(n_1807), .ZN(n_1600));
   INV_X1 i_367 (.A(n_1602), .ZN(n_1601));
   OAI22_X1 i_368 (.A1(n_1745), .A2(n_1746), .B1(n_1808), .B2(n_1604), .ZN(
      n_1602));
   OAI21_X1 i_369 (.A(n_1809), .B1(n_1745), .B2(n_1746), .ZN(n_1603));
   OAI21_X1 i_370 (.A(n_1792), .B1(n_1800), .B2(n_1605), .ZN(n_1604));
   INV_X1 i_371 (.A(n_1606), .ZN(n_1605));
   OAI21_X1 i_372 (.A(n_1797), .B1(n_1803), .B2(n_1607), .ZN(n_1606));
   INV_X1 i_373 (.A(n_893), .ZN(n_1607));
   OAI22_X1 i_374 (.A1(n_1742), .A2(n_1739), .B1(n_1820), .B2(n_1821), .ZN(
      n_1609));
   XOR2_X1 i_375 (.A(n_1782), .B(n_1616), .Z(mult_res[33]));
   XOR2_X1 i_376 (.A(n_1780), .B(n_1612), .Z(mult_res[34]));
   XNOR2_X1 i_377 (.A(n_1617), .B(n_1611), .ZN(mult_res[36]));
   OAI22_X1 i_378 (.A1(n_1735), .A2(n_1771), .B1(n_1775), .B2(n_1778), .ZN(
      n_1611));
   AOI21_X1 i_379 (.A(n_1815), .B1(n_1733), .B2(n_1734), .ZN(n_1612));
   OAI21_X1 i_380 (.A(n_1781), .B1(n_1740), .B2(n_1732), .ZN(n_1616));
   NOR2_X1 i_381 (.A1(n_1680), .A2(n_1671), .ZN(n_1617));
   XOR2_X1 i_382 (.A(n_1667), .B(n_1624), .Z(mult_res[37]));
   XOR2_X1 i_383 (.A(n_1623), .B(n_1620), .Z(mult_res[38]));
   XOR2_X1 i_384 (.A(n_1621), .B(n_1618), .Z(mult_res[39]));
   NOR2_X1 i_385 (.A1(n_1664), .A2(n_1655), .ZN(n_1618));
   XNOR2_X1 i_386 (.A(n_1625), .B(n_1619), .ZN(mult_res[40]));
   OAI22_X1 i_387 (.A1(n_955), .A2(n_968), .B1(n_1655), .B2(n_1621), .ZN(n_1619));
   AOI21_X1 i_388 (.A(n_1665), .B1(n_939), .B2(n_954), .ZN(n_1620));
   AOI21_X1 i_389 (.A(n_1665), .B1(n_1659), .B2(n_1622), .ZN(n_1621));
   INV_X1 i_390 (.A(n_1623), .ZN(n_1622));
   AOI21_X1 i_391 (.A(n_1662), .B1(n_1667), .B2(n_1660), .ZN(n_1623));
   OAI21_X1 i_392 (.A(n_1660), .B1(n_921), .B2(n_938), .ZN(n_1624));
   NOR2_X1 i_393 (.A1(n_1666), .A2(n_1657), .ZN(n_1625));
   XOR2_X1 i_394 (.A(n_1653), .B(n_1632), .Z(mult_res[41]));
   XOR2_X1 i_395 (.A(n_1631), .B(n_1630), .Z(mult_res[42]));
   XNOR2_X1 i_396 (.A(n_1627), .B(n_1626), .ZN(mult_res[43]));
   OAI22_X1 i_397 (.A1(n_991), .A2(n_998), .B1(n_1643), .B2(n_1631), .ZN(n_1626));
   NOR2_X1 i_398 (.A1(n_1650), .A2(n_1639), .ZN(n_1627));
   XNOR2_X1 i_399 (.A(n_1633), .B(n_1628), .ZN(mult_res[44]));
   OAI22_X1 i_400 (.A1(n_1631), .A2(n_1629), .B1(n_1649), .B2(n_1639), .ZN(
      n_1628));
   NAND2_X1 i_401 (.A1(n_1640), .A2(n_1630), .ZN(n_1629));
   NOR2_X1 i_402 (.A1(n_1651), .A2(n_1643), .ZN(n_1630));
   AOI21_X1 i_403 (.A(n_1647), .B1(n_1653), .B2(n_1645), .ZN(n_1631));
   OAI21_X1 i_404 (.A(n_1645), .B1(n_981), .B2(n_990), .ZN(n_1632));
   NOR2_X1 i_405 (.A1(n_1652), .A2(n_1641), .ZN(n_1633));
   XOR2_X1 i_406 (.A(n_1637), .B(n_1634), .Z(mult_res[45]));
   AOI21_X1 i_407 (.A(n_1763), .B1(n_1768), .B2(n_1767), .ZN(n_1634));
   XNOR2_X1 i_408 (.A(n_1636), .B(n_1635), .ZN(mult_res[46]));
   AOI21_X1 i_409 (.A(n_1765), .B1(n_1011), .B2(n_1766), .ZN(n_1635));
   AOI21_X1 i_410 (.A(n_1765), .B1(n_1764), .B2(n_1636), .ZN(mult_res[47]));
   OAI22_X1 i_411 (.A1(n_1009), .A2(n_1010), .B1(n_1763), .B2(n_1637), .ZN(
      n_1636));
   OR4_X1 i_412 (.A1(n_1641), .A2(n_1638), .A3(n_1642), .A4(n_1646), .ZN(n_1637));
   NOR2_X1 i_413 (.A1(n_1652), .A2(n_1640), .ZN(n_1638));
   INV_X1 i_414 (.A(n_1640), .ZN(n_1639));
   NAND2_X1 i_415 (.A1(n_999), .A2(n_1004), .ZN(n_1640));
   AND2_X1 i_416 (.A1(n_1005), .A2(n_1008), .ZN(n_1641));
   AOI21_X1 i_417 (.A(n_1648), .B1(n_1645), .B2(n_1644), .ZN(n_1642));
   INV_X1 i_418 (.A(n_1644), .ZN(n_1643));
   NAND2_X1 i_419 (.A1(n_991), .A2(n_998), .ZN(n_1644));
   NAND2_X1 i_420 (.A1(n_981), .A2(n_990), .ZN(n_1645));
   NOR3_X1 i_421 (.A1(n_1648), .A2(n_1647), .A3(n_1653), .ZN(n_1646));
   NOR2_X1 i_422 (.A1(n_981), .A2(n_990), .ZN(n_1647));
   OAI21_X1 i_423 (.A(n_1649), .B1(n_1005), .B2(n_1008), .ZN(n_1648));
   NOR2_X1 i_424 (.A1(n_1651), .A2(n_1650), .ZN(n_1649));
   NOR2_X1 i_425 (.A1(n_999), .A2(n_1004), .ZN(n_1650));
   NOR2_X1 i_426 (.A1(n_991), .A2(n_998), .ZN(n_1651));
   NOR2_X1 i_427 (.A1(n_1005), .A2(n_1008), .ZN(n_1652));
   NOR4_X1 i_428 (.A1(n_1657), .A2(n_1654), .A3(n_1658), .A4(n_1661), .ZN(n_1653));
   NOR2_X1 i_429 (.A1(n_1666), .A2(n_1656), .ZN(n_1654));
   INV_X1 i_430 (.A(n_1656), .ZN(n_1655));
   NAND2_X1 i_431 (.A1(n_955), .A2(n_968), .ZN(n_1656));
   AND2_X1 i_432 (.A1(n_969), .A2(n_980), .ZN(n_1657));
   AOI21_X1 i_433 (.A(n_1663), .B1(n_1660), .B2(n_1659), .ZN(n_1658));
   NAND2_X1 i_434 (.A1(n_939), .A2(n_954), .ZN(n_1659));
   NAND2_X1 i_435 (.A1(n_921), .A2(n_938), .ZN(n_1660));
   NOR3_X1 i_436 (.A1(n_1663), .A2(n_1662), .A3(n_1667), .ZN(n_1661));
   NOR2_X1 i_437 (.A1(n_921), .A2(n_938), .ZN(n_1662));
   OR3_X1 i_438 (.A1(n_1666), .A2(n_1664), .A3(n_1665), .ZN(n_1663));
   NOR2_X1 i_439 (.A1(n_955), .A2(n_968), .ZN(n_1664));
   NOR2_X1 i_440 (.A1(n_939), .A2(n_954), .ZN(n_1665));
   NOR2_X1 i_441 (.A1(n_969), .A2(n_980), .ZN(n_1666));
   NOR4_X1 i_442 (.A1(n_1671), .A2(n_1668), .A3(n_1672), .A4(n_1675), .ZN(n_1667));
   NOR2_X1 i_443 (.A1(n_1680), .A2(n_1776), .ZN(n_1668));
   AND2_X1 i_444 (.A1(n_1772), .A2(n_920), .ZN(n_1671));
   AOI21_X1 i_445 (.A(n_1677), .B1(n_1781), .B2(n_1814), .ZN(n_1672));
   NOR3_X1 i_446 (.A1(n_1677), .A2(n_1813), .A3(n_1782), .ZN(n_1675));
   OR3_X1 i_447 (.A1(n_1680), .A2(n_1777), .A3(n_1815), .ZN(n_1677));
   NOR2_X1 i_448 (.A1(n_1772), .A2(n_920), .ZN(n_1680));
   OAI222_X1 i_449 (.A1(n_881), .A2(n_883), .B1(n_2), .B2(n_4), .C1(n_1695), 
      .C2(n_1692), .ZN(n_659));
   AOI211_X1 i_450 (.A(n_1701), .B(n_1693), .C1(n_1670), .C2(n_1773), .ZN(n_1692));
   AOI22_X1 i_451 (.A1(Na[2]), .A2(n_0), .B1(Na[0]), .B2(n_1694), .ZN(n_1693));
   NOR2_X1 i_452 (.A1(n_1702), .A2(n_1669), .ZN(n_1694));
   AND2_X1 i_453 (.A1(n_2), .A2(n_4), .ZN(n_1695));
   INV_X1 i_454 (.A(n_1795), .ZN(n_1717));
   NOR2_X1 i_455 (.A1(n_1750), .A2(n_1753), .ZN(n_668));
   NOR2_X1 i_456 (.A1(n_1748), .A2(n_1749), .ZN(n_669));
   NOR2_X1 i_457 (.A1(n_1754), .A2(n_1744), .ZN(n_670));
   NOR2_X1 i_458 (.A1(n_1768), .A2(n_1767), .ZN(n_1763));
   NAND2_X1 i_459 (.A1(n_1011), .A2(n_1766), .ZN(n_1764));
   NOR2_X1 i_460 (.A1(n_1011), .A2(n_1766), .ZN(n_1765));
   NOR2_X1 i_461 (.A1(n_1725), .A2(n_1700), .ZN(n_1766));
   INV_X1 i_462 (.A(n_1010), .ZN(n_1767));
   INV_X1 i_463 (.A(n_1009), .ZN(n_1768));
   INV_X1 i_464 (.A(n_0), .ZN(n_1773));
   FA_X1 i_465 (.A(n_1451), .B(n_1474), .CI(n_1497), .CO(n_353), .S(n_352));
   FA_X1 i_466 (.A(n_1382), .B(n_1405), .CI(n_1428), .CO(n_351), .S(n_350));
   FA_X1 i_467 (.A(n_1313), .B(n_1336), .CI(n_1359), .CO(n_349), .S(n_348));
   FA_X1 i_468 (.A(n_352), .B(n_350), .CI(n_348), .CO(n_363), .S(n_362));
   FA_X1 i_469 (.A(n_1430), .B(n_1453), .CI(n_1476), .CO(n_281), .S(n_280));
   FA_X1 i_470 (.A(n_1361), .B(n_1384), .CI(n_1407), .CO(n_279), .S(n_278));
   FA_X1 i_471 (.A(n_1292), .B(n_1315), .CI(n_1338), .CO(n_277), .S(n_276));
   FA_X1 i_472 (.A(n_281), .B(n_279), .CI(n_277), .CO(n_321), .S(n_320));
   FA_X1 i_473 (.A(n_1499), .B(n_1522), .CI(n_1545), .CO(n_283), .S(n_282));
   FA_X1 i_474 (.A(n_1544), .B(n_1565), .CI(n_283), .CO(n_319), .S(n_318));
   FA_X1 i_475 (.A(n_1520), .B(n_1543), .CI(n_1564), .CO(n_355), .S(n_354));
   FA_X1 i_476 (.A(n_321), .B(n_319), .CI(n_354), .CO(n_361), .S(n_360));
   FA_X1 i_477 (.A(n_1223), .B(n_1246), .CI(n_1269), .CO(n_275), .S(n_274));
   FA_X1 i_478 (.A(n_1154), .B(n_1177), .CI(n_1200), .CO(n_273), .S(n_272));
   FA_X1 i_479 (.A(n_1385), .B(n_1408), .CI(n_1431), .CO(n_247), .S(n_246));
   FA_X1 i_480 (.A(n_1316), .B(n_1339), .CI(n_1362), .CO(n_245), .S(n_244));
   FA_X1 i_481 (.A(n_1247), .B(n_1270), .CI(n_1293), .CO(n_243), .S(n_242));
   FA_X1 i_482 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_287), .S(n_286));
   FA_X1 i_483 (.A(n_275), .B(n_273), .CI(n_287), .CO(n_323), .S(n_322));
   FA_X1 i_484 (.A(n_1268), .B(n_1291), .CI(n_1314), .CO(n_311), .S(n_310));
   FA_X1 i_485 (.A(n_1199), .B(n_1222), .CI(n_1245), .CO(n_309), .S(n_308));
   FA_X1 i_486 (.A(n_1130), .B(n_1153), .CI(n_1176), .CO(n_307), .S(n_306));
   FA_X1 i_487 (.A(n_311), .B(n_309), .CI(n_307), .CO(n_359), .S(n_358));
   FA_X1 i_488 (.A(n_1475), .B(n_1498), .CI(n_1521), .CO(n_317), .S(n_316));
   FA_X1 i_489 (.A(n_1406), .B(n_1429), .CI(n_1452), .CO(n_315), .S(n_314));
   FA_X1 i_490 (.A(n_1337), .B(n_1360), .CI(n_1383), .CO(n_313), .S(n_312));
   FA_X1 i_491 (.A(n_317), .B(n_315), .CI(n_313), .CO(n_357), .S(n_356));
   FA_X1 i_492 (.A(n_323), .B(n_358), .CI(n_356), .CO(n_367), .S(n_366));
   FA_X1 i_493 (.A(n_363), .B(n_361), .CI(n_367), .CO(n_409), .S(n_408));
   FA_X1 i_494 (.A(n_1427), .B(n_1450), .CI(n_1473), .CO(n_391), .S(n_390));
   FA_X1 i_495 (.A(n_1358), .B(n_1381), .CI(n_1404), .CO(n_389), .S(n_388));
   FA_X1 i_496 (.A(n_1289), .B(n_1312), .CI(n_1335), .CO(n_387), .S(n_386));
   FA_X1 i_497 (.A(n_391), .B(n_389), .CI(n_387), .CO(n_437), .S(n_436));
   FA_X1 i_498 (.A(n_1220), .B(n_1243), .CI(n_1266), .CO(n_385), .S(n_384));
   FA_X1 i_499 (.A(n_388), .B(n_386), .CI(n_384), .CO(n_403), .S(n_402));
   FA_X1 i_500 (.A(n_1496), .B(n_1519), .CI(n_1542), .CO(n_393), .S(n_392));
   FA_X1 i_501 (.A(n_357), .B(n_392), .CI(n_390), .CO(n_401), .S(n_400));
   FA_X1 i_502 (.A(n_436), .B(n_403), .CI(n_401), .CO(n_449), .S(n_448));
   FA_X1 i_503 (.A(n_1151), .B(n_1174), .CI(n_1197), .CO(n_383), .S(n_382));
   FA_X1 i_504 (.A(n_1082), .B(n_1105), .CI(n_1128), .CO(n_381), .S(n_380));
   FA_X1 i_505 (.A(n_1175), .B(n_1198), .CI(n_1221), .CO(n_345), .S(n_344));
   FA_X1 i_506 (.A(n_1106), .B(n_1129), .CI(n_1152), .CO(n_343), .S(n_342));
   FA_X1 i_507 (.A(n_345), .B(n_343), .CI(n_359), .CO(n_399), .S(n_398));
   FA_X1 i_508 (.A(n_382), .B(n_380), .CI(n_398), .CO(n_405), .S(n_404));
   FA_X1 i_509 (.A(n_404), .B(n_402), .CI(n_400), .CO(n_411), .S(n_410));
   FA_X1 i_510 (.A(n_409), .B(n_448), .CI(n_411), .CO(n_455), .S(n_454));
   FA_X1 i_511 (.A(n_280), .B(n_278), .CI(n_276), .CO(n_291), .S(n_290));
   FA_X1 i_512 (.A(n_1178), .B(n_1201), .CI(n_1224), .CO(n_241), .S(n_240));
   FA_X1 i_513 (.A(n_1478), .B(n_1501), .CI(n_1524), .CO(n_219), .S(n_218));
   FA_X1 i_514 (.A(n_1409), .B(n_1432), .CI(n_1455), .CO(n_217), .S(n_216));
   FA_X1 i_515 (.A(n_1340), .B(n_1363), .CI(n_1386), .CO(n_215), .S(n_214));
   FA_X1 i_516 (.A(n_219), .B(n_217), .CI(n_215), .CO(n_253), .S(n_252));
   FA_X1 i_517 (.A(n_241), .B(n_253), .CI(n_282), .CO(n_289), .S(n_288));
   FA_X1 i_518 (.A(n_320), .B(n_291), .CI(n_289), .CO(n_331), .S(n_330));
   FA_X1 i_519 (.A(n_308), .B(n_306), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_520 (.A(n_1244), .B(n_1267), .CI(n_1290), .CO(n_347), .S(n_346));
   FA_X1 i_521 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_365), .S(n_364));
   FA_X1 i_522 (.A(n_331), .B(n_329), .CI(n_364), .CO(n_371), .S(n_370));
   FA_X1 i_523 (.A(n_314), .B(n_312), .CI(n_310), .CO(n_327), .S(n_326));
   FA_X1 i_524 (.A(n_1523), .B(n_1546), .CI(n_1567), .CO(n_251), .S(n_250));
   FA_X1 i_525 (.A(n_1454), .B(n_1477), .CI(n_1500), .CO(n_249), .S(n_248));
   FA_X1 i_526 (.A(n_1566), .B(n_251), .CI(n_249), .CO(n_285), .S(n_284));
   FA_X1 i_527 (.A(n_285), .B(n_318), .CI(n_316), .CO(n_325), .S(n_324));
   FA_X1 i_528 (.A(n_327), .B(n_325), .CI(n_360), .CO(n_369), .S(n_368));
   FA_X1 i_529 (.A(n_362), .B(n_368), .CI(n_366), .CO(n_373), .S(n_372));
   FA_X1 i_530 (.A(n_371), .B(n_373), .CI(n_410), .CO(n_415), .S(n_414));
   FA_X1 i_531 (.A(n_351), .B(n_349), .CI(n_347), .CO(n_397), .S(n_396));
   FA_X1 i_532 (.A(n_1563), .B(n_355), .CI(n_353), .CO(n_395), .S(n_394));
   FA_X1 i_533 (.A(n_1541), .B(n_1562), .CI(n_393), .CO(n_435), .S(n_434));
   FA_X1 i_534 (.A(n_397), .B(n_395), .CI(n_434), .CO(n_441), .S(n_440));
   FA_X1 i_535 (.A(n_396), .B(n_394), .CI(n_365), .CO(n_407), .S(n_406));
   FA_X1 i_536 (.A(n_440), .B(n_407), .CI(n_405), .CO(n_451), .S(n_450));
   FA_X1 i_537 (.A(n_369), .B(n_408), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_538 (.A(n_1265), .B(n_1288), .CI(n_1311), .CO(n_427), .S(n_426));
   FA_X1 i_539 (.A(n_1196), .B(n_1219), .CI(n_1242), .CO(n_425), .S(n_424));
   FA_X1 i_540 (.A(n_1127), .B(n_1150), .CI(n_1173), .CO(n_423), .S(n_422));
   FA_X1 i_541 (.A(n_426), .B(n_424), .CI(n_422), .CO(n_445), .S(n_444));
   FA_X1 i_542 (.A(n_1472), .B(n_1495), .CI(n_1518), .CO(n_433), .S(n_432));
   FA_X1 i_543 (.A(n_1403), .B(n_1426), .CI(n_1449), .CO(n_431), .S(n_430));
   FA_X1 i_544 (.A(n_1334), .B(n_1357), .CI(n_1380), .CO(n_429), .S(n_428));
   FA_X1 i_545 (.A(n_432), .B(n_430), .CI(n_428), .CO(n_443), .S(n_442));
   FA_X1 i_546 (.A(n_1058), .B(n_1081), .CI(n_1104), .CO(n_421), .S(n_420));
   FA_X1 i_547 (.A(n_385), .B(n_383), .CI(n_381), .CO(n_439), .S(n_438));
   FA_X1 i_548 (.A(n_420), .B(n_399), .CI(n_438), .CO(n_447), .S(n_446));
   FA_X1 i_549 (.A(n_444), .B(n_442), .CI(n_446), .CO(n_453), .S(n_452));
   FA_X1 i_550 (.A(n_450), .B(n_413), .CI(n_452), .CO(n_457), .S(n_456));
   FA_X1 i_551 (.A(n_454), .B(n_415), .CI(n_456), .CO(n_459), .S(n_458));
   FA_X1 i_552 (.A(n_421), .B(n_439), .CI(n_437), .CO(n_483), .S(n_482));
   FA_X1 i_553 (.A(n_443), .B(n_441), .CI(n_482), .CO(n_493), .S(n_492));
   FA_X1 i_554 (.A(n_427), .B(n_425), .CI(n_423), .CO(n_481), .S(n_480));
   FA_X1 i_555 (.A(n_433), .B(n_431), .CI(n_429), .CO(n_479), .S(n_478));
   FA_X1 i_556 (.A(n_480), .B(n_478), .CI(n_445), .CO(n_491), .S(n_490));
   FA_X1 i_557 (.A(n_492), .B(n_490), .CI(n_453), .CO(n_499), .S(n_498));
   FA_X1 i_558 (.A(n_1172), .B(n_1195), .CI(n_1218), .CO(n_467), .S(n_466));
   FA_X1 i_559 (.A(n_1103), .B(n_1126), .CI(n_1149), .CO(n_465), .S(n_464));
   FA_X1 i_560 (.A(n_1034), .B(n_1057), .CI(n_1080), .CO(n_463), .S(n_462));
   FA_X1 i_561 (.A(n_466), .B(n_464), .CI(n_462), .CO(n_489), .S(n_488));
   FA_X1 i_562 (.A(n_449), .B(n_447), .CI(n_488), .CO(n_495), .S(n_494));
   FA_X1 i_563 (.A(n_1379), .B(n_1402), .CI(n_1425), .CO(n_473), .S(n_472));
   FA_X1 i_564 (.A(n_1310), .B(n_1333), .CI(n_1356), .CO(n_471), .S(n_470));
   FA_X1 i_565 (.A(n_1241), .B(n_1264), .CI(n_1287), .CO(n_469), .S(n_468));
   FA_X1 i_566 (.A(n_472), .B(n_470), .CI(n_468), .CO(n_487), .S(n_486));
   FA_X1 i_567 (.A(n_1517), .B(n_1540), .CI(n_1561), .CO(n_477), .S(n_476));
   FA_X1 i_568 (.A(n_1448), .B(n_1471), .CI(n_1494), .CO(n_475), .S(n_474));
   FA_X1 i_569 (.A(n_435), .B(n_476), .CI(n_474), .CO(n_485), .S(n_484));
   FA_X1 i_570 (.A(n_486), .B(n_484), .CI(n_451), .CO(n_497), .S(n_496));
   FA_X1 i_571 (.A(n_494), .B(n_455), .CI(n_496), .CO(n_501), .S(n_500));
   FA_X1 i_572 (.A(n_498), .B(n_457), .CI(n_500), .CO(n_503), .S(n_502));
   HA_X1 i_573 (.A(n_459), .B(n_502), .CO(n_684), .S(n_682));
   FA_X1 i_574 (.A(n_469), .B(n_467), .CI(n_465), .CO(n_686), .S(n_524));
   FA_X1 i_575 (.A(n_475), .B(n_473), .CI(n_471), .CO(n_688), .S(n_522));
   FA_X1 i_576 (.A(n_524), .B(n_522), .CI(n_489), .CO(n_690), .S(n_534));
   FA_X1 i_577 (.A(n_534), .B(n_495), .CI(n_497), .CO(n_692), .S(n_542));
   FA_X1 i_578 (.A(n_1102), .B(n_1125), .CI(n_1148), .CO(n_694), .S(n_508));
   FA_X1 i_579 (.A(n_1033), .B(n_1056), .CI(n_1079), .CO(n_696), .S(n_506));
   FA_X1 i_580 (.A(n_508), .B(n_506), .CI(n_483), .CO(n_697), .S(n_532));
   FA_X1 i_581 (.A(n_1309), .B(n_1332), .CI(n_1355), .CO(n_698), .S(n_514));
   FA_X1 i_582 (.A(n_1240), .B(n_1263), .CI(n_1286), .CO(n_699), .S(n_512));
   FA_X1 i_583 (.A(n_1171), .B(n_1194), .CI(n_1217), .CO(n_704), .S(n_510));
   FA_X1 i_584 (.A(n_514), .B(n_512), .CI(n_510), .CO(n_705), .S(n_530));
   FA_X1 i_585 (.A(n_491), .B(n_532), .CI(n_530), .CO(n_724), .S(n_538));
   FA_X1 i_586 (.A(n_1516), .B(n_1539), .CI(n_477), .CO(n_726), .S(n_520));
   FA_X1 i_587 (.A(n_1447), .B(n_1470), .CI(n_1493), .CO(n_732), .S(n_518));
   FA_X1 i_588 (.A(n_1378), .B(n_1401), .CI(n_1424), .CO(n_733), .S(n_516));
   FA_X1 i_589 (.A(n_520), .B(n_518), .CI(n_516), .CO(n_738), .S(n_528));
   FA_X1 i_590 (.A(n_463), .B(n_481), .CI(n_479), .CO(n_771), .S(n_526));
   FA_X1 i_591 (.A(n_487), .B(n_485), .CI(n_526), .CO(n_800), .S(n_536));
   FA_X1 i_592 (.A(n_528), .B(n_493), .CI(n_536), .CO(n_801), .S(n_540));
   FA_X1 i_593 (.A(n_499), .B(n_538), .CI(n_540), .CO(n_828), .S(n_544));
   FA_X1 i_594 (.A(n_542), .B(n_501), .CI(n_544), .CO(n_829), .S(n_546));
   HA_X1 i_595 (.A(n_503), .B(n_546), .CO(n_855), .S(n_854));
   FA_X1 i_596 (.A(n_1271), .B(n_1294), .CI(n_1317), .CO(n_213), .S(n_212));
   FA_X1 i_597 (.A(n_1202), .B(n_1225), .CI(n_1248), .CO(n_211), .S(n_210));
   FA_X1 i_598 (.A(n_1433), .B(n_1456), .CI(n_1479), .CO(n_189), .S(n_188));
   FA_X1 i_599 (.A(n_1364), .B(n_1387), .CI(n_1410), .CO(n_187), .S(n_186));
   FA_X1 i_600 (.A(n_1295), .B(n_1318), .CI(n_1341), .CO(n_185), .S(n_184));
   FA_X1 i_601 (.A(n_189), .B(n_187), .CI(n_185), .CO(n_223), .S(n_222));
   FA_X1 i_602 (.A(n_213), .B(n_211), .CI(n_223), .CO(n_255), .S(n_254));
   FA_X1 i_603 (.A(n_274), .B(n_272), .CI(n_255), .CO(n_293), .S(n_292));
   FA_X1 i_604 (.A(n_246), .B(n_244), .CI(n_242), .CO(n_259), .S(n_258));
   FA_X1 i_605 (.A(n_286), .B(n_284), .CI(n_259), .CO(n_295), .S(n_294));
   FA_X1 i_606 (.A(n_293), .B(n_295), .CI(n_328), .CO(n_333), .S(n_332));
   FA_X1 i_607 (.A(n_1502), .B(n_1525), .CI(n_1548), .CO(n_191), .S(n_190));
   FA_X1 i_608 (.A(n_1547), .B(n_1568), .CI(n_191), .CO(n_221), .S(n_220));
   FA_X1 i_609 (.A(n_221), .B(n_250), .CI(n_248), .CO(n_257), .S(n_256));
   FA_X1 i_610 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_229), .S(n_228));
   FA_X1 i_611 (.A(n_220), .B(n_218), .CI(n_216), .CO(n_227), .S(n_226));
   FA_X1 i_612 (.A(n_252), .B(n_229), .CI(n_227), .CO(n_263), .S(n_262));
   FA_X1 i_613 (.A(n_257), .B(n_288), .CI(n_263), .CO(n_297), .S(n_296));
   FA_X1 i_614 (.A(n_326), .B(n_324), .CI(n_297), .CO(n_335), .S(n_334));
   FA_X1 i_615 (.A(n_333), .B(n_335), .CI(n_370), .CO(n_375), .S(n_374));
   FA_X1 i_616 (.A(n_375), .B(n_412), .CI(n_414), .CO(n_417), .S(n_416));
   HA_X1 i_617 (.A(n_417), .B(n_458), .CO(n_878), .S(n_460));
   FA_X1 i_618 (.A(n_595), .B(n_597), .CI(n_599), .CO(n_183), .S(n_182));
   FA_X1 i_619 (.A(n_158), .B(n_156), .CI(n_140), .CO(n_195), .S(n_194));
   FA_X1 i_620 (.A(n_657), .B(n_162), .CI(n_160), .CO(n_193), .S(n_192));
   FA_X1 i_621 (.A(n_183), .B(n_195), .CI(n_193), .CO(n_225), .S(n_224));
   FA_X1 i_622 (.A(n_240), .B(n_225), .CI(n_254), .CO(n_261), .S(n_260));
   FA_X1 i_623 (.A(n_261), .B(n_292), .CI(n_290), .CO(n_299), .S(n_298));
   FA_X1 i_624 (.A(n_330), .B(n_299), .CI(n_332), .CO(n_337), .S(n_336));
   FA_X1 i_625 (.A(n_337), .B(n_372), .CI(n_374), .CO(n_377), .S(n_376));
   HA_X1 i_626 (.A(n_377), .B(n_416), .CO(n_419), .S(n_418));
   FA_X1 i_627 (.A(n_222), .B(n_199), .CI(n_197), .CO(n_231), .S(n_230));
   FA_X1 i_628 (.A(n_231), .B(n_258), .CI(n_256), .CO(n_265), .S(n_264));
   FA_X1 i_629 (.A(n_294), .B(n_265), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_630 (.A(n_334), .B(n_301), .CI(n_336), .CO(n_339), .S(n_338));
   FA_X1 i_631 (.A(n_224), .B(n_201), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_632 (.A(n_260), .B(n_262), .CI(n_233), .CO(n_267), .S(n_266));
   FA_X1 i_633 (.A(n_267), .B(n_298), .CI(n_300), .CO(n_303), .S(n_302));
   HA_X1 i_634 (.A(n_303), .B(n_338), .CO(n_341), .S(n_340));
   HA_X1 i_635 (.A(n_339), .B(n_341), .CO(n_379), .S(n_378));
   FA_X1 i_636 (.A(n_226), .B(n_230), .CI(n_203), .CO(n_235), .S(n_234));
   FA_X1 i_637 (.A(n_235), .B(n_264), .CI(n_266), .CO(n_269), .S(n_268));
   HA_X1 i_638 (.A(n_269), .B(n_302), .CO(n_305), .S(n_304));
   FA_X1 i_639 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_640 (.A(n_232), .B(n_205), .CI(n_234), .CO(n_237), .S(n_236));
   FA_X1 i_641 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_642 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   HA_X1 i_643 (.A(n_207), .B(n_209), .CO(n_239), .S(n_238));
   HA_X1 i_644 (.A(n_237), .B(n_239), .CO(n_271), .S(n_270));
   FA_X1 i_645 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_646 (.A(n_143), .B(n_138), .CI(n_163), .CO(n_173), .S(n_172));
   FA_X1 i_647 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_171), .S(n_170));
   FA_X1 i_648 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_649 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_650 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_651 (.A(n_164), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_652 (.A(n_147), .B(n_145), .CI(n_165), .CO(n_175), .S(n_174));
   FA_X1 i_653 (.A(n_166), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_654 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_655 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   FA_X1 i_656 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_657 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   HA_X1 i_658 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_659 (.A(n_91), .B(n_85), .CI(n_96), .CO(n_121), .S(n_120));
   FA_X1 i_660 (.A(n_113), .B(n_111), .CI(n_99), .CO(n_879), .S(n_142));
   FA_X1 i_661 (.A(n_114), .B(n_112), .CI(n_110), .CO(n_123), .S(n_122));
   FA_X1 i_662 (.A(n_66), .B(n_93), .CI(n_92), .CO(n_101), .S(n_100));
   FA_X1 i_663 (.A(n_90), .B(n_84), .CI(n_67), .CO(n_103), .S(n_102));
   FA_X1 i_664 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_665 (.A(n_94), .B(n_81), .CI(n_83), .CO(n_105), .S(n_104));
   FA_X1 i_666 (.A(n_98), .B(n_120), .CI(n_115), .CO(n_125), .S(n_124));
   FA_X1 i_667 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   FA_X1 i_668 (.A(n_132), .B(n_119), .CI(n_118), .CO(n_147), .S(n_146));
   FA_X1 i_669 (.A(n_116), .B(n_136), .CI(n_134), .CO(n_145), .S(n_144));
   FA_X1 i_670 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_671 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   HA_X1 i_672 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_673 (.A(n_64), .B(n_79), .CI(n_82), .CO(n_87), .S(n_86));
   HA_X1 i_674 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_675 (.A(n_48), .B(n_50), .CI(n_51), .CO(n_69), .S(n_68));
   HA_X1 i_676 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_677 (.A(n_24), .B(n_22), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_678 (.A(n_30), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_679 (.A(n_36), .B(n_32), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_680 (.A(n_39), .B(n_37), .CO(n_55), .S(n_54));
   FA_X1 i_681 (.A(n_14), .B(n_12), .CI(n_20), .CO(n_27), .S(n_26));
   HA_X1 i_682 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_683 (.A(n_7), .B(n_8), .CI(n_10), .CO(n_17), .S(n_16));
   HA_X1 i_684 (.A(n_9), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_685 (.A(n_609), .B(n_630), .CI(n_631), .CO(n_7), .S(n_881));
   HA_X1 i_686 (.A(n_3), .B(n_6), .CO(n_11), .S(n_883));
   NOR2_X1 i_687 (.A1(n_1702), .A2(n_1687), .ZN(n_1548));
   NOR2_X1 i_688 (.A1(n_1703), .A2(n_1686), .ZN(n_1525));
   NOR2_X1 i_689 (.A1(n_1704), .A2(n_1685), .ZN(n_1502));
   NOR2_X1 i_690 (.A1(n_1701), .A2(n_1689), .ZN(n_1568));
   NOR2_X1 i_691 (.A1(n_1702), .A2(n_1688), .ZN(n_1547));
   NOR2_X1 i_692 (.A1(n_1711), .A2(n_1676), .ZN(n_1341));
   NOR2_X1 i_693 (.A1(n_1712), .A2(n_1674), .ZN(n_1318));
   NOR2_X1 i_694 (.A1(n_1713), .A2(n_1673), .ZN(n_1295));
   NOR2_X1 i_695 (.A1(n_1708), .A2(n_1681), .ZN(n_1410));
   NOR2_X1 i_696 (.A1(n_1709), .A2(n_1679), .ZN(n_1387));
   NOR2_X1 i_697 (.A1(n_1710), .A2(n_1678), .ZN(n_1364));
   NOR2_X1 i_698 (.A1(n_1705), .A2(n_1684), .ZN(n_1479));
   NOR2_X1 i_699 (.A1(n_1706), .A2(n_1683), .ZN(n_1456));
   NOR2_X1 i_700 (.A1(n_1707), .A2(n_1682), .ZN(n_1433));
   NOR2_X1 i_701 (.A1(n_1715), .A2(n_1670), .ZN(n_1248));
   NOR2_X1 i_702 (.A1(n_1716), .A2(n_1669), .ZN(n_1225));
   NOR2_X1 i_703 (.A1(n_1718), .A2(n_1615), .ZN(n_1202));
   NOR2_X1 i_704 (.A1(n_1712), .A2(n_1676), .ZN(n_1317));
   NOR2_X1 i_705 (.A1(n_1713), .A2(n_1674), .ZN(n_1294));
   NOR2_X1 i_706 (.A1(n_1714), .A2(n_1673), .ZN(n_1271));
   NOR2_X1 i_707 (.A1(n_1707), .A2(n_1691), .ZN(n_1424));
   NOR2_X1 i_708 (.A1(n_1708), .A2(n_1690), .ZN(n_1401));
   NOR2_X1 i_709 (.A1(n_1709), .A2(n_1689), .ZN(n_1378));
   NOR2_X1 i_710 (.A1(n_1704), .A2(n_1698), .ZN(n_1493));
   NOR2_X1 i_711 (.A1(n_1705), .A2(n_1697), .ZN(n_1470));
   NOR2_X1 i_712 (.A1(n_1706), .A2(n_1696), .ZN(n_1447));
   NOR2_X1 i_713 (.A1(n_1702), .A2(n_1700), .ZN(n_1539));
   NOR2_X1 i_714 (.A1(n_1703), .A2(n_1699), .ZN(n_1516));
   NOR2_X1 i_715 (.A1(n_1716), .A2(n_1682), .ZN(n_1217));
   NOR2_X1 i_716 (.A1(n_1718), .A2(n_1681), .ZN(n_1194));
   NOR2_X1 i_717 (.A1(n_1719), .A2(n_1679), .ZN(n_1171));
   NOR2_X1 i_718 (.A1(n_1713), .A2(n_1685), .ZN(n_1286));
   NOR2_X1 i_719 (.A1(n_1714), .A2(n_1684), .ZN(n_1263));
   NOR2_X1 i_720 (.A1(n_1715), .A2(n_1683), .ZN(n_1240));
   NOR2_X1 i_721 (.A1(n_1710), .A2(n_1688), .ZN(n_1355));
   NOR2_X1 i_722 (.A1(n_1711), .A2(n_1687), .ZN(n_1332));
   NOR2_X1 i_723 (.A1(n_1712), .A2(n_1686), .ZN(n_1309));
   NOR2_X1 i_724 (.A1(n_1723), .A2(n_1673), .ZN(n_1079));
   NOR2_X1 i_725 (.A1(n_1724), .A2(n_1670), .ZN(n_1056));
   NOR2_X1 i_726 (.A1(n_1725), .A2(n_1669), .ZN(n_1033));
   NOR2_X1 i_727 (.A1(n_1720), .A2(n_1678), .ZN(n_1148));
   NOR2_X1 i_728 (.A1(n_1721), .A2(n_1676), .ZN(n_1125));
   NOR2_X1 i_729 (.A1(n_1722), .A2(n_1674), .ZN(n_1102));
   NOR2_X1 i_730 (.A1(n_1704), .A2(n_1697), .ZN(n_1494));
   NOR2_X1 i_731 (.A1(n_1705), .A2(n_1696), .ZN(n_1471));
   NOR2_X1 i_732 (.A1(n_1706), .A2(n_1691), .ZN(n_1448));
   NOR2_X1 i_733 (.A1(n_1701), .A2(n_1700), .ZN(n_1561));
   NOR2_X1 i_734 (.A1(n_1702), .A2(n_1699), .ZN(n_1540));
   NOR2_X1 i_735 (.A1(n_1703), .A2(n_1698), .ZN(n_1517));
   NOR2_X1 i_736 (.A1(n_1713), .A2(n_1684), .ZN(n_1287));
   NOR2_X1 i_737 (.A1(n_1714), .A2(n_1683), .ZN(n_1264));
   NOR2_X1 i_738 (.A1(n_1715), .A2(n_1682), .ZN(n_1241));
   NOR2_X1 i_739 (.A1(n_1710), .A2(n_1687), .ZN(n_1356));
   NOR2_X1 i_740 (.A1(n_1711), .A2(n_1686), .ZN(n_1333));
   NOR2_X1 i_741 (.A1(n_1712), .A2(n_1685), .ZN(n_1310));
   NOR2_X1 i_742 (.A1(n_1707), .A2(n_1690), .ZN(n_1425));
   NOR2_X1 i_743 (.A1(n_1708), .A2(n_1689), .ZN(n_1402));
   NOR2_X1 i_745 (.A1(n_1709), .A2(n_1688), .ZN(n_1379));
   NOR2_X1 i_746 (.A1(n_1723), .A2(n_1670), .ZN(n_1080));
   NOR2_X1 i_747 (.A1(n_1724), .A2(n_1669), .ZN(n_1057));
   NOR2_X1 i_748 (.A1(n_1725), .A2(n_1615), .ZN(n_1034));
   NOR2_X1 i_749 (.A1(n_1720), .A2(n_1676), .ZN(n_1149));
   NOR2_X1 i_750 (.A1(n_1721), .A2(n_1674), .ZN(n_1126));
   NOR2_X1 i_751 (.A1(n_1722), .A2(n_1673), .ZN(n_1103));
   NOR2_X1 i_752 (.A1(n_1716), .A2(n_1681), .ZN(n_1218));
   NOR2_X1 i_753 (.A1(n_1718), .A2(n_1679), .ZN(n_1195));
   NOR2_X1 i_754 (.A1(n_1719), .A2(n_1678), .ZN(n_1172));
   NOR2_X1 i_755 (.A1(n_1722), .A2(n_1670), .ZN(n_1104));
   NOR2_X1 i_756 (.A1(n_1723), .A2(n_1669), .ZN(n_1081));
   NOR2_X1 i_757 (.A1(n_1724), .A2(n_1615), .ZN(n_1058));
   NOR2_X1 i_758 (.A1(n_1709), .A2(n_1687), .ZN(n_1380));
   NOR2_X1 i_759 (.A1(n_1710), .A2(n_1686), .ZN(n_1357));
   NOR2_X1 i_760 (.A1(n_1711), .A2(n_1685), .ZN(n_1334));
   NOR2_X1 i_761 (.A1(n_1706), .A2(n_1690), .ZN(n_1449));
   NOR2_X1 i_762 (.A1(n_1707), .A2(n_1689), .ZN(n_1426));
   NOR2_X1 i_763 (.A1(n_1708), .A2(n_1688), .ZN(n_1403));
   NOR2_X1 i_764 (.A1(n_1703), .A2(n_1697), .ZN(n_1518));
   NOR2_X1 i_765 (.A1(n_1704), .A2(n_1696), .ZN(n_1495));
   NOR2_X1 i_766 (.A1(n_1705), .A2(n_1691), .ZN(n_1472));
   NOR2_X1 i_768 (.A1(n_1719), .A2(n_1676), .ZN(n_1173));
   NOR2_X1 i_769 (.A1(n_1720), .A2(n_1674), .ZN(n_1150));
   NOR2_X1 i_770 (.A1(n_1721), .A2(n_1673), .ZN(n_1127));
   NOR2_X1 i_771 (.A1(n_1715), .A2(n_1681), .ZN(n_1242));
   NOR2_X1 i_772 (.A1(n_1716), .A2(n_1679), .ZN(n_1219));
   NOR2_X1 i_773 (.A1(n_1718), .A2(n_1678), .ZN(n_1196));
   NOR2_X1 i_774 (.A1(n_1712), .A2(n_1684), .ZN(n_1311));
   NOR2_X1 i_775 (.A1(n_1713), .A2(n_1683), .ZN(n_1288));
   NOR2_X1 i_776 (.A1(n_1714), .A2(n_1682), .ZN(n_1265));
   NOR2_X1 i_777 (.A1(n_1701), .A2(n_1699), .ZN(n_1562));
   NOR2_X1 i_778 (.A1(n_1702), .A2(n_1698), .ZN(n_1541));
   NOR2_X1 i_779 (.A1(n_1701), .A2(n_1698), .ZN(n_1563));
   NOR2_X1 i_780 (.A1(n_1704), .A2(n_1687), .ZN(n_1500));
   NOR2_X1 i_781 (.A1(n_1705), .A2(n_1686), .ZN(n_1477));
   NOR2_X1 i_782 (.A1(n_1706), .A2(n_1685), .ZN(n_1454));
   NOR2_X1 i_783 (.A1(n_1701), .A2(n_1690), .ZN(n_1567));
   NOR2_X1 i_784 (.A1(n_1702), .A2(n_1689), .ZN(n_1546));
   NOR2_X1 i_785 (.A1(n_1703), .A2(n_1688), .ZN(n_1523));
   NOR2_X1 i_786 (.A1(n_1701), .A2(n_1691), .ZN(n_1566));
   NOR2_X1 i_787 (.A1(n_1713), .A2(n_1681), .ZN(n_1290));
   NOR2_X1 i_788 (.A1(n_1714), .A2(n_1679), .ZN(n_1267));
   NOR2_X1 i_789 (.A1(n_1715), .A2(n_1678), .ZN(n_1244));
   NOR2_X1 i_791 (.A1(n_1709), .A2(n_1681), .ZN(n_1386));
   NOR2_X1 i_793 (.A1(n_1710), .A2(n_1679), .ZN(n_1363));
   NOR2_X1 i_794 (.A1(n_1711), .A2(n_1678), .ZN(n_1340));
   NOR2_X1 i_795 (.A1(n_1706), .A2(n_1684), .ZN(n_1455));
   NOR2_X1 i_796 (.A1(n_1707), .A2(n_1683), .ZN(n_1432));
   NOR2_X1 i_797 (.A1(n_1708), .A2(n_1682), .ZN(n_1409));
   NOR2_X1 i_798 (.A1(n_1703), .A2(n_1687), .ZN(n_1524));
   NOR2_X1 i_799 (.A1(n_1704), .A2(n_1686), .ZN(n_1501));
   NOR2_X1 i_800 (.A1(n_1705), .A2(n_1685), .ZN(n_1478));
   NOR2_X1 i_801 (.A1(n_1716), .A2(n_1670), .ZN(n_1224));
   NOR2_X1 i_802 (.A1(n_1718), .A2(n_1669), .ZN(n_1201));
   NOR2_X1 i_803 (.A1(n_1719), .A2(n_1615), .ZN(n_1178));
   NOR2_X1 i_804 (.A1(n_1720), .A2(n_1670), .ZN(n_1152));
   NOR2_X1 i_805 (.A1(n_1721), .A2(n_1669), .ZN(n_1129));
   NOR2_X1 i_806 (.A1(n_1722), .A2(n_1615), .ZN(n_1106));
   NOR2_X1 i_807 (.A1(n_1716), .A2(n_1676), .ZN(n_1221));
   NOR2_X1 i_808 (.A1(n_1718), .A2(n_1674), .ZN(n_1198));
   NOR2_X1 i_809 (.A1(n_1719), .A2(n_1673), .ZN(n_1175));
   NOR2_X1 i_810 (.A1(n_1721), .A2(n_1670), .ZN(n_1128));
   NOR2_X1 i_811 (.A1(n_1722), .A2(n_1669), .ZN(n_1105));
   NOR2_X1 i_812 (.A1(n_1723), .A2(n_1615), .ZN(n_1082));
   NOR2_X1 i_814 (.A1(n_1718), .A2(n_1676), .ZN(n_1197));
   NOR2_X1 i_817 (.A1(n_1719), .A2(n_1674), .ZN(n_1174));
   NOR2_X1 i_818 (.A1(n_1720), .A2(n_1673), .ZN(n_1151));
   NOR2_X1 i_819 (.A1(n_1702), .A2(n_1697), .ZN(n_1542));
   NOR2_X1 i_820 (.A1(n_1703), .A2(n_1696), .ZN(n_1519));
   NOR2_X1 i_821 (.A1(n_1704), .A2(n_1691), .ZN(n_1496));
   NOR2_X1 i_822 (.A1(n_1714), .A2(n_1681), .ZN(n_1266));
   NOR2_X1 i_823 (.A1(n_1715), .A2(n_1679), .ZN(n_1243));
   NOR2_X1 i_824 (.A1(n_1716), .A2(n_1678), .ZN(n_1220));
   NOR2_X1 i_825 (.A1(n_1711), .A2(n_1684), .ZN(n_1335));
   NOR2_X1 i_826 (.A1(n_1712), .A2(n_1683), .ZN(n_1312));
   NOR2_X1 i_827 (.A1(n_1713), .A2(n_1682), .ZN(n_1289));
   NOR2_X1 i_828 (.A1(n_1708), .A2(n_1687), .ZN(n_1404));
   NOR2_X1 i_829 (.A1(n_1709), .A2(n_1686), .ZN(n_1381));
   NOR2_X1 i_830 (.A1(n_1710), .A2(n_1685), .ZN(n_1358));
   NOR2_X1 i_831 (.A1(n_1705), .A2(n_1690), .ZN(n_1473));
   NOR2_X1 i_832 (.A1(n_1706), .A2(n_1689), .ZN(n_1450));
   NOR2_X1 i_833 (.A1(n_1707), .A2(n_1688), .ZN(n_1427));
   NOR2_X1 i_834 (.A1(n_1709), .A2(n_1684), .ZN(n_1383));
   NOR2_X1 i_835 (.A1(n_1710), .A2(n_1683), .ZN(n_1360));
   NOR2_X1 i_837 (.A1(n_1711), .A2(n_1682), .ZN(n_1337));
   NOR2_X1 i_840 (.A1(n_1706), .A2(n_1687), .ZN(n_1452));
   NOR2_X1 i_841 (.A1(n_1707), .A2(n_1686), .ZN(n_1429));
   NOR2_X1 i_842 (.A1(n_1708), .A2(n_1685), .ZN(n_1406));
   NOR2_X1 i_843 (.A1(n_1703), .A2(n_1690), .ZN(n_1521));
   NOR2_X1 i_844 (.A1(n_1704), .A2(n_1689), .ZN(n_1498));
   NOR2_X1 i_845 (.A1(n_1705), .A2(n_1688), .ZN(n_1475));
   NOR2_X1 i_846 (.A1(n_1719), .A2(n_1670), .ZN(n_1176));
   NOR2_X1 i_847 (.A1(n_1720), .A2(n_1669), .ZN(n_1153));
   NOR2_X1 i_848 (.A1(n_1721), .A2(n_1615), .ZN(n_1130));
   NOR2_X1 i_849 (.A1(n_1715), .A2(n_1676), .ZN(n_1245));
   NOR2_X1 i_850 (.A1(n_1716), .A2(n_1674), .ZN(n_1222));
   NOR2_X1 i_851 (.A1(n_1718), .A2(n_1673), .ZN(n_1199));
   NOR2_X1 i_852 (.A1(n_1712), .A2(n_1681), .ZN(n_1314));
   NOR2_X1 i_853 (.A1(n_1713), .A2(n_1679), .ZN(n_1291));
   NOR2_X1 i_854 (.A1(n_1714), .A2(n_1678), .ZN(n_1268));
   NOR2_X1 i_855 (.A1(n_1713), .A2(n_1676), .ZN(n_1293));
   NOR2_X1 i_856 (.A1(n_1714), .A2(n_1674), .ZN(n_1270));
   NOR2_X1 i_857 (.A1(n_1715), .A2(n_1673), .ZN(n_1247));
   NOR2_X1 i_858 (.A1(n_1710), .A2(n_1681), .ZN(n_1362));
   NOR2_X1 i_860 (.A1(n_1711), .A2(n_1679), .ZN(n_1339));
   NOR2_X1 i_863 (.A1(n_1712), .A2(n_1678), .ZN(n_1316));
   NOR2_X1 i_864 (.A1(n_1707), .A2(n_1684), .ZN(n_1431));
   NOR2_X1 i_865 (.A1(n_1708), .A2(n_1683), .ZN(n_1408));
   NOR2_X1 i_866 (.A1(n_1709), .A2(n_1682), .ZN(n_1385));
   NOR2_X1 i_867 (.A1(n_1718), .A2(n_1670), .ZN(n_1200));
   NOR2_X1 i_868 (.A1(n_1719), .A2(n_1669), .ZN(n_1177));
   NOR2_X1 i_869 (.A1(n_1720), .A2(n_1615), .ZN(n_1154));
   NOR2_X1 i_870 (.A1(n_1714), .A2(n_1676), .ZN(n_1269));
   NOR2_X1 i_871 (.A1(n_1715), .A2(n_1674), .ZN(n_1246));
   NOR2_X1 i_872 (.A1(n_1716), .A2(n_1673), .ZN(n_1223));
   NOR2_X1 i_873 (.A1(n_1701), .A2(n_1697), .ZN(n_1564));
   NOR2_X1 i_874 (.A1(n_1702), .A2(n_1696), .ZN(n_1543));
   NOR2_X1 i_875 (.A1(n_1703), .A2(n_1691), .ZN(n_1520));
   NOR2_X1 i_876 (.A1(n_1702), .A2(n_1690), .ZN(n_1545));
   NOR2_X1 i_877 (.A1(n_1703), .A2(n_1689), .ZN(n_1522));
   NOR2_X1 i_878 (.A1(n_1704), .A2(n_1688), .ZN(n_1499));
   NOR2_X1 i_879 (.A1(n_1701), .A2(n_1696), .ZN(n_1565));
   NOR2_X1 i_880 (.A1(n_1702), .A2(n_1691), .ZN(n_1544));
   NOR2_X1 i_881 (.A1(n_1711), .A2(n_1681), .ZN(n_1338));
   NOR2_X1 i_883 (.A1(n_1712), .A2(n_1679), .ZN(n_1315));
   NOR2_X1 i_886 (.A1(n_1713), .A2(n_1678), .ZN(n_1292));
   NOR2_X1 i_887 (.A1(n_1708), .A2(n_1684), .ZN(n_1407));
   NOR2_X1 i_888 (.A1(n_1709), .A2(n_1683), .ZN(n_1384));
   NOR2_X1 i_889 (.A1(n_1710), .A2(n_1682), .ZN(n_1361));
   NOR2_X1 i_890 (.A1(n_1705), .A2(n_1687), .ZN(n_1476));
   NOR2_X1 i_891 (.A1(n_1706), .A2(n_1686), .ZN(n_1453));
   NOR2_X1 i_892 (.A1(n_1707), .A2(n_1685), .ZN(n_1430));
   NOR2_X1 i_893 (.A1(n_1710), .A2(n_1684), .ZN(n_1359));
   NOR2_X1 i_894 (.A1(n_1711), .A2(n_1683), .ZN(n_1336));
   NOR2_X1 i_895 (.A1(n_1712), .A2(n_1682), .ZN(n_1313));
   NOR2_X1 i_896 (.A1(n_1707), .A2(n_1687), .ZN(n_1428));
   NOR2_X1 i_897 (.A1(n_1708), .A2(n_1686), .ZN(n_1405));
   NOR2_X1 i_898 (.A1(n_1709), .A2(n_1685), .ZN(n_1382));
   NOR2_X1 i_899 (.A1(n_1704), .A2(n_1690), .ZN(n_1497));
   NOR2_X1 i_900 (.A1(n_1705), .A2(n_1689), .ZN(n_1474));
   NOR2_X1 i_901 (.A1(n_1706), .A2(n_1688), .ZN(n_1451));
   XNOR2_X1 i_902 (.A(n_887), .B(n_885), .ZN(mult_res[24]));
   OAI22_X1 i_903 (.A1(n_682), .A2(n_878), .B1(n_1583), .B2(n_889), .ZN(n_885));
   AOI21_X1 i_904 (.A(n_1585), .B1(n_684), .B2(n_854), .ZN(n_887));
   AOI21_X1 i_906 (.A(n_1569), .B1(n_1536), .B2(n_891), .ZN(n_889));
   OAI21_X1 i_909 (.A(n_1513), .B1(n_1490), .B2(n_893), .ZN(n_891));
   NAND2_X1 i_910 (.A1(n_1329), .A2(n_895), .ZN(n_893));
   OAI211_X1 i_911 (.A(n_897), .B(n_1421), .C1(n_268), .C2(n_270), .ZN(n_895));
   OAI221_X1 i_912 (.A(n_901), .B1(n_1053), .B2(n_900), .C1(n_1076), .C2(n_899), 
      .ZN(n_897));
   AOI22_X1 i_913 (.A1(n_236), .A2(n_238), .B1(n_206), .B2(n_208), .ZN(n_899));
   AOI22_X1 i_914 (.A1(n_152), .A2(n_154), .B1(n_178), .B2(n_180), .ZN(n_900));
   OAI211_X1 i_915 (.A(n_1030), .B(n_1099), .C1(n_152), .C2(n_154), .ZN(n_901));
   INV_X1 i_916 (.A(n_1053), .ZN(n_1030));
   OAI222_X1 i_917 (.A1(n_178), .A2(n_180), .B1(n_206), .B2(n_208), .C1(n_236), 
      .C2(n_238), .ZN(n_1053));
   NOR2_X1 i_918 (.A1(n_236), .A2(n_238), .ZN(n_1076));
   OAI211_X1 i_919 (.A(n_1145), .B(n_1122), .C1(n_1226), .C2(n_1168), .ZN(n_1099));
   AOI21_X1 i_920 (.A(n_1191), .B1(n_128), .B2(n_130), .ZN(n_1122));
   OAI211_X1 i_921 (.A(n_106), .B(n_108), .C1(n_128), .C2(n_130), .ZN(n_1145));
   AOI22_X1 i_922 (.A1(n_68), .A2(n_70), .B1(n_86), .B2(n_88), .ZN(n_1168));
   AOI211_X1 i_923 (.A(n_1226), .B(n_1214), .C1(n_1306), .C2(n_1237), .ZN(n_1191));
   OAI22_X1 i_924 (.A1(n_68), .A2(n_70), .B1(n_52), .B2(n_54), .ZN(n_1214));
   OAI222_X1 i_925 (.A1(n_86), .A2(n_88), .B1(n_106), .B2(n_108), .C1(n_128), 
      .C2(n_130), .ZN(n_1226));
   OAI221_X1 i_926 (.A(n_1249), .B1(n_26), .B2(n_28), .C1(n_38), .C2(n_40), 
      .ZN(n_1237));
   OAI21_X1 i_927 (.A(n_1283), .B1(n_1272), .B2(n_1260), .ZN(n_1249));
   NOR2_X1 i_929 (.A1(n_16), .A2(n_18), .ZN(n_1260));
   AOI21_X1 i_932 (.A(n_1614), .B1(n_881), .B2(n_883), .ZN(n_1272));
   AOI22_X1 i_933 (.A1(n_16), .A2(n_18), .B1(n_26), .B2(n_28), .ZN(n_1283));
   AOI22_X1 i_934 (.A1(n_52), .A2(n_54), .B1(n_38), .B2(n_40), .ZN(n_1306));
   AOI221_X1 i_935 (.A(n_1352), .B1(n_1421), .B2(n_1375), .C1(n_376), .C2(n_378), 
      .ZN(n_1329));
   NOR3_X1 i_936 (.A1(n_1610), .A2(n_1444), .A3(n_1586), .ZN(n_1352));
   INV_X1 i_937 (.A(n_1398), .ZN(n_1375));
   AOI22_X1 i_938 (.A1(n_268), .A2(n_270), .B1(n_304), .B2(n_271), .ZN(n_1398));
   AOI211_X1 i_939 (.A(n_1444), .B(n_1467), .C1(n_1610), .C2(n_1586), .ZN(n_1421));
   NOR2_X1 i_940 (.A1(n_376), .A2(n_378), .ZN(n_1444));
   NOR2_X1 i_941 (.A1(n_304), .A2(n_271), .ZN(n_1467));
   NOR2_X1 i_942 (.A1(n_1613), .A2(n_1608), .ZN(n_1490));
   NAND2_X1 i_943 (.A1(n_1613), .A2(n_1608), .ZN(n_1513));
   NAND2_X1 i_944 (.A1(n_460), .A2(n_419), .ZN(n_1536));
   NOR2_X1 i_945 (.A1(n_460), .A2(n_419), .ZN(n_1569));
   INV_X1 i_946 (.A(n_1584), .ZN(n_1583));
   NAND2_X1 i_947 (.A1(n_682), .A2(n_878), .ZN(n_1584));
   NOR2_X1 i_948 (.A1(n_684), .A2(n_854), .ZN(n_1585));
   INV_X1 i_949 (.A(n_305), .ZN(n_1586));
   INV_X1 i_950 (.A(n_379), .ZN(n_1608));
   INV_X1 i_952 (.A(n_340), .ZN(n_1610));
   INV_X1 i_955 (.A(n_418), .ZN(n_1613));
   INV_X1 i_956 (.A(n_659), .ZN(n_1614));
   INV_X1 i_957 (.A(Na[0]), .ZN(n_1615));
   INV_X1 i_958 (.A(Na[1]), .ZN(n_1669));
   INV_X1 i_959 (.A(Na[2]), .ZN(n_1670));
   INV_X1 i_960 (.A(Na[3]), .ZN(n_1673));
   INV_X1 i_961 (.A(Na[4]), .ZN(n_1674));
   INV_X1 i_962 (.A(Na[5]), .ZN(n_1676));
   INV_X1 i_963 (.A(Na[6]), .ZN(n_1678));
   INV_X1 i_964 (.A(Na[7]), .ZN(n_1679));
   INV_X1 i_965 (.A(Na[8]), .ZN(n_1681));
   INV_X1 i_966 (.A(Na[9]), .ZN(n_1682));
   INV_X1 i_967 (.A(Na[10]), .ZN(n_1683));
   INV_X1 i_968 (.A(Na[11]), .ZN(n_1684));
   INV_X1 i_969 (.A(Na[12]), .ZN(n_1685));
   INV_X1 i_970 (.A(Na[13]), .ZN(n_1686));
   INV_X1 i_971 (.A(Na[14]), .ZN(n_1687));
   INV_X1 i_972 (.A(Na[15]), .ZN(n_1688));
   INV_X1 i_973 (.A(Na[16]), .ZN(n_1689));
   INV_X1 i_975 (.A(Na[17]), .ZN(n_1690));
   INV_X1 i_978 (.A(Na[18]), .ZN(n_1691));
   INV_X1 i_979 (.A(Na[19]), .ZN(n_1696));
   INV_X1 i_980 (.A(Na[20]), .ZN(n_1697));
   INV_X1 i_981 (.A(Na[21]), .ZN(n_1698));
   INV_X1 i_982 (.A(Na[22]), .ZN(n_1699));
   INV_X1 i_983 (.A(Na[23]), .ZN(n_1700));
   INV_X1 i_984 (.A(Nb[0]), .ZN(n_1701));
   INV_X1 i_985 (.A(Nb[1]), .ZN(n_1702));
   INV_X1 i_986 (.A(Nb[2]), .ZN(n_1703));
   INV_X1 i_987 (.A(Nb[3]), .ZN(n_1704));
   INV_X1 i_988 (.A(Nb[4]), .ZN(n_1705));
   INV_X1 i_989 (.A(Nb[5]), .ZN(n_1706));
   INV_X1 i_990 (.A(Nb[6]), .ZN(n_1707));
   INV_X1 i_991 (.A(Nb[7]), .ZN(n_1708));
   INV_X1 i_992 (.A(Nb[8]), .ZN(n_1709));
   INV_X1 i_993 (.A(Nb[9]), .ZN(n_1710));
   INV_X1 i_994 (.A(Nb[10]), .ZN(n_1711));
   INV_X1 i_995 (.A(Nb[11]), .ZN(n_1712));
   INV_X1 i_996 (.A(Nb[12]), .ZN(n_1713));
   INV_X1 i_998 (.A(Nb[13]), .ZN(n_1714));
   INV_X1 i_999 (.A(Nb[14]), .ZN(n_1715));
   INV_X1 i_1001 (.A(Nb[15]), .ZN(n_1716));
   INV_X1 i_1002 (.A(Nb[16]), .ZN(n_1718));
   INV_X1 i_1003 (.A(Nb[17]), .ZN(n_1719));
   INV_X1 i_1004 (.A(Nb[18]), .ZN(n_1720));
   INV_X1 i_1005 (.A(Nb[19]), .ZN(n_1721));
   INV_X1 i_1006 (.A(Nb[20]), .ZN(n_1722));
   INV_X1 i_1007 (.A(Nb[21]), .ZN(n_1723));
   INV_X1 i_1008 (.A(Nb[22]), .ZN(n_1724));
   INV_X1 i_1009 (.A(Nb[23]), .ZN(n_1725));
   FA_X1 i_1010 (.A(n_1095), .B(n_1118), .CI(n_1141), .CO(n_775), .S(n_774));
   FA_X1 i_1011 (.A(n_1026), .B(n_1049), .CI(n_1072), .CO(n_773), .S(n_772));
   FA_X1 i_1012 (.A(n_1165), .B(n_1188), .CI(n_1211), .CO(n_745), .S(n_744));
   FA_X1 i_1013 (.A(n_1096), .B(n_1119), .CI(n_1142), .CO(n_743), .S(n_742));
   FA_X1 i_1014 (.A(n_1027), .B(n_1050), .CI(n_1073), .CO(n_741), .S(n_740));
   FA_X1 i_1015 (.A(n_745), .B(n_743), .CI(n_741), .CO(n_785), .S(n_784));
   FA_X1 i_1016 (.A(n_775), .B(n_773), .CI(n_785), .CO(n_815), .S(n_814));
   FA_X1 i_1017 (.A(n_1302), .B(n_1325), .CI(n_1348), .CO(n_781), .S(n_780));
   FA_X1 i_1018 (.A(n_1233), .B(n_1256), .CI(n_1279), .CO(n_779), .S(n_778));
   FA_X1 i_1019 (.A(n_1164), .B(n_1187), .CI(n_1210), .CO(n_777), .S(n_776));
   FA_X1 i_1021 (.A(n_781), .B(n_779), .CI(n_777), .CO(n_813), .S(n_812));
   FA_X1 i_1022 (.A(n_778), .B(n_776), .CI(n_774), .CO(n_789), .S(n_788));
   FA_X1 i_1024 (.A(n_814), .B(n_812), .CI(n_789), .CO(n_821), .S(n_820));
   FA_X1 i_1025 (.A(n_1231), .B(n_1254), .CI(n_1277), .CO(n_837), .S(n_836));
   FA_X1 i_1026 (.A(n_1162), .B(n_1185), .CI(n_1208), .CO(n_835), .S(n_834));
   FA_X1 i_1027 (.A(n_1093), .B(n_1116), .CI(n_1139), .CO(n_833), .S(n_832));
   FA_X1 i_1028 (.A(n_836), .B(n_834), .CI(n_832), .CO(n_845), .S(n_844));
   FA_X1 i_1029 (.A(n_1024), .B(n_1047), .CI(n_1070), .CO(n_831), .S(n_830));
   FA_X1 i_1030 (.A(n_1232), .B(n_1255), .CI(n_1278), .CO(n_809), .S(n_808));
   FA_X1 i_1031 (.A(n_1163), .B(n_1186), .CI(n_1209), .CO(n_807), .S(n_806));
   FA_X1 i_1032 (.A(n_1094), .B(n_1117), .CI(n_1140), .CO(n_805), .S(n_804));
   FA_X1 i_1033 (.A(n_809), .B(n_807), .CI(n_805), .CO(n_841), .S(n_840));
   FA_X1 i_1034 (.A(n_830), .B(n_815), .CI(n_840), .CO(n_847), .S(n_846));
   FA_X1 i_1035 (.A(n_821), .B(n_844), .CI(n_846), .CO(n_851), .S(n_850));
   FA_X1 i_1036 (.A(n_1304), .B(n_1327), .CI(n_1350), .CO(n_715), .S(n_714));
   FA_X1 i_1037 (.A(n_1235), .B(n_1258), .CI(n_1281), .CO(n_713), .S(n_712));
   FA_X1 i_1038 (.A(n_1166), .B(n_1189), .CI(n_1212), .CO(n_711), .S(n_710));
   FA_X1 i_1039 (.A(n_715), .B(n_713), .CI(n_711), .CO(n_753), .S(n_752));
   FA_X1 i_1040 (.A(n_1373), .B(n_1396), .CI(n_1419), .CO(n_717), .S(n_716));
   FA_X1 i_1041 (.A(n_1372), .B(n_1395), .CI(n_717), .CO(n_751), .S(n_750));
   FA_X1 i_1042 (.A(n_753), .B(n_751), .CI(n_780), .CO(n_787), .S(n_786));
   FA_X1 i_1044 (.A(n_1303), .B(n_1326), .CI(n_1349), .CO(n_749), .S(n_748));
   FA_X1 i_1045 (.A(n_1234), .B(n_1257), .CI(n_1280), .CO(n_747), .S(n_746));
   FA_X1 i_1047 (.A(n_1371), .B(n_749), .CI(n_747), .CO(n_783), .S(n_782));
   FA_X1 i_1048 (.A(n_746), .B(n_744), .CI(n_742), .CO(n_759), .S(n_758));
   FA_X1 i_1049 (.A(n_1374), .B(n_1397), .CI(n_1420), .CO(n_681), .S(n_680));
   FA_X1 i_1050 (.A(n_1305), .B(n_1328), .CI(n_1351), .CO(n_679), .S(n_678));
   FA_X1 i_1051 (.A(n_1236), .B(n_1259), .CI(n_1282), .CO(n_677), .S(n_676));
   FA_X1 i_1052 (.A(n_681), .B(n_679), .CI(n_677), .CO(n_719), .S(n_718));
   FA_X1 i_1054 (.A(n_719), .B(n_750), .CI(n_748), .CO(n_757), .S(n_756));
   FA_X1 i_1055 (.A(n_782), .B(n_759), .CI(n_757), .CO(n_793), .S(n_792));
   FA_X1 i_1056 (.A(n_1097), .B(n_1120), .CI(n_1143), .CO(n_709), .S(n_708));
   FA_X1 i_1057 (.A(n_1028), .B(n_1051), .CI(n_1074), .CO(n_707), .S(n_706));
   FA_X1 i_1058 (.A(n_1167), .B(n_1190), .CI(n_1213), .CO(n_675), .S(n_674));
   FA_X1 i_1059 (.A(n_1098), .B(n_1121), .CI(n_1144), .CO(n_673), .S(n_672));
   FA_X1 i_1060 (.A(n_1029), .B(n_1052), .CI(n_1075), .CO(n_671), .S(n_1726));
   FA_X1 i_1061 (.A(n_675), .B(n_673), .CI(n_671), .CO(n_721), .S(n_720));
   FA_X1 i_1062 (.A(n_709), .B(n_707), .CI(n_721), .CO(n_755), .S(n_754));
   FA_X1 i_1063 (.A(n_772), .B(n_755), .CI(n_784), .CO(n_791), .S(n_790));
   FA_X1 i_1065 (.A(n_787), .B(n_793), .CI(n_791), .CO(n_823), .S(n_822));
   FA_X1 i_1068 (.A(n_788), .B(n_790), .CI(n_792), .CO(n_797), .S(n_796));
   FA_X1 i_1069 (.A(n_820), .B(n_822), .CI(n_797), .CO(n_827), .S(n_826));
   FA_X1 i_1070 (.A(n_1025), .B(n_1048), .CI(n_1071), .CO(n_803), .S(n_802));
   FA_X1 i_1071 (.A(n_806), .B(n_804), .CI(n_802), .CO(n_819), .S(n_818));
   FA_X1 i_1072 (.A(n_1301), .B(n_1324), .CI(n_1347), .CO(n_811), .S(n_810));
   FA_X1 i_1073 (.A(n_783), .B(n_810), .CI(n_808), .CO(n_817), .S(n_816));
   FA_X1 i_1075 (.A(n_1300), .B(n_1323), .CI(n_811), .CO(n_839), .S(n_838));
   FA_X1 i_1076 (.A(n_803), .B(n_813), .CI(n_838), .CO(n_843), .S(n_842));
   FA_X1 i_1077 (.A(n_819), .B(n_817), .CI(n_842), .CO(n_849), .S(n_848));
   FA_X1 i_1078 (.A(n_740), .B(n_754), .CI(n_752), .CO(n_761), .S(n_760));
   FA_X1 i_1079 (.A(n_714), .B(n_712), .CI(n_710), .CO(n_725), .S(n_1727));
   FA_X1 i_1080 (.A(n_596), .B(n_598), .CI(n_600), .CO(n_639), .S(n_638));
   FA_X1 i_1081 (.A(n_592), .B(n_593), .CI(n_594), .CO(n_637), .S(n_636));
   FA_X1 i_1082 (.A(n_579), .B(n_590), .CI(n_591), .CO(n_635), .S(n_634));
   FA_X1 i_1083 (.A(n_639), .B(n_637), .CI(n_635), .CO(n_685), .S(n_1728));
   FA_X1 i_1084 (.A(n_604), .B(n_605), .CI(n_606), .CO(n_643), .S(n_642));
   FA_X1 i_1085 (.A(n_601), .B(n_602), .CI(n_603), .CO(n_641), .S(n_640));
   FA_X1 i_1086 (.A(n_1443), .B(n_643), .CI(n_641), .CO(n_683), .S(n_1729));
   FA_X1 i_1087 (.A(n_685), .B(n_683), .CI(n_716), .CO(n_723), .S(n_722));
   FA_X1 i_1088 (.A(n_574), .B(n_575), .CI(n_578), .CO(n_633), .S(n_632));
   FA_X1 i_1089 (.A(n_533), .B(n_529), .CI(n_525), .CO(n_649), .S(n_648));
   FA_X1 i_1090 (.A(n_545), .B(n_541), .CI(n_537), .CO(n_647), .S(n_646));
   FA_X1 i_1091 (.A(n_633), .B(n_649), .CI(n_647), .CO(n_687), .S(n_1730));
   FA_X1 i_1092 (.A(n_708), .B(n_706), .CI(n_687), .CO(n_727), .S(n_1731));
   FA_X1 i_1093 (.A(n_725), .B(n_723), .CI(n_727), .CO(n_763), .S(n_762));
   FA_X1 i_1094 (.A(n_786), .B(n_761), .CI(n_763), .CO(n_795), .S(n_794));
   FA_X1 i_1095 (.A(n_818), .B(n_816), .CI(n_795), .CO(n_825), .S(n_824));
   FA_X1 i_1096 (.A(n_823), .B(n_848), .CI(n_825), .CO(n_853), .S(n_852));
   FA_X1 i_1097 (.A(n_850), .B(n_827), .CI(n_852), .CO(n_1733), .S(n_1732));
   FA_X1 i_1098 (.A(n_1092), .B(n_1115), .CI(n_1138), .CO(n_859), .S(n_858));
   FA_X1 i_1099 (.A(n_1023), .B(n_1046), .CI(n_1069), .CO(n_857), .S(n_856));
   FA_X1 i_1100 (.A(n_833), .B(n_831), .CI(n_841), .CO(n_867), .S(n_866));
   FA_X1 i_1101 (.A(n_858), .B(n_856), .CI(n_866), .CO(n_871), .S(n_870));
   FA_X1 i_1102 (.A(n_1230), .B(n_1253), .CI(n_1276), .CO(n_863), .S(n_862));
   FA_X1 i_1103 (.A(n_1161), .B(n_1184), .CI(n_1207), .CO(n_861), .S(n_860));
   FA_X1 i_1104 (.A(n_839), .B(n_862), .CI(n_860), .CO(n_869), .S(n_868));
   FA_X1 i_1105 (.A(n_847), .B(n_870), .CI(n_868), .CO(n_875), .S(n_874));
   FA_X1 i_1106 (.A(n_1299), .B(n_837), .CI(n_835), .CO(n_865), .S(n_864));
   FA_X1 i_1107 (.A(n_864), .B(n_845), .CI(n_843), .CO(n_873), .S(n_872));
   FA_X1 i_1108 (.A(n_849), .B(n_872), .CI(n_851), .CO(n_877), .S(n_876));
   FA_X1 i_1109 (.A(n_853), .B(n_874), .CI(n_876), .CO(n_1735), .S(n_1734));
   FA_X1 i_1110 (.A(n_676), .B(n_674), .CI(n_672), .CO(n_691), .S(n_1736));
   FA_X1 i_1111 (.A(n_720), .B(n_718), .CI(n_691), .CO(n_729), .S(n_728));
   FA_X1 i_1112 (.A(n_729), .B(n_758), .CI(n_756), .CO(n_765), .S(n_764));
   FA_X1 i_1113 (.A(n_607), .B(n_608), .CI(n_548), .CO(n_645), .S(n_644));
   FA_X1 i_1114 (.A(n_645), .B(n_680), .CI(n_678), .CO(n_689), .S(n_1737));
   FA_X1 i_1115 (.A(n_636), .B(n_634), .CI(n_632), .CO(n_655), .S(n_654));
   FA_X1 i_1116 (.A(n_642), .B(n_640), .CI(n_638), .CO(n_653), .S(n_652));
   FA_X1 i_1117 (.A(n_566), .B(n_551), .CI(n_644), .CO(n_651), .S(n_650));
   FA_X1 i_1118 (.A(n_655), .B(n_653), .CI(n_651), .CO(n_695), .S(n_1738));
   FA_X1 i_1119 (.A(n_689), .B(n_722), .CI(n_695), .CO(n_731), .S(n_730));
   FA_X1 i_1120 (.A(n_731), .B(n_762), .CI(n_760), .CO(n_767), .S(n_766));
   FA_X1 i_1121 (.A(n_765), .B(n_794), .CI(n_767), .CO(n_799), .S(n_798));
   FA_X1 i_1122 (.A(n_824), .B(n_799), .CI(n_826), .CO(n_1740), .S(n_1739));
   FA_X1 i_1123 (.A(n_573), .B(n_764), .CI(n_735), .CO(n_769), .S(n_768));
   FA_X1 i_1124 (.A(n_796), .B(n_769), .CI(n_798), .CO(n_1742), .S(n_1741));
   FA_X1 i_1125 (.A(n_571), .B(n_572), .CI(n_701), .CO(n_737), .S(n_736));
   FA_X1 i_1126 (.A(n_766), .B(n_737), .CI(n_768), .CO(n_1743), .S(n_770));
   FA_X1 i_1127 (.A(n_567), .B(n_661), .CI(n_568), .CO(n_701), .S(n_700));
   FA_X1 i_1128 (.A(n_625), .B(n_662), .CI(n_627), .CO(n_667), .S(n_666));
   FA_X1 i_1129 (.A(n_663), .B(n_570), .CI(n_665), .CO(n_703), .S(n_702));
   FA_X1 i_1130 (.A(n_700), .B(n_667), .CI(n_702), .CO(n_1745), .S(n_1744));
   FA_X1 i_1131 (.A(n_728), .B(n_569), .CI(n_730), .CO(n_735), .S(n_734));
   FA_X1 i_1132 (.A(n_734), .B(n_703), .CI(n_736), .CO(n_739), .S(n_1746));
   FA_X1 i_1133 (.A(n_586), .B(n_588), .CI(n_829), .CO(n_1748), .S(n_1747));
   FA_X1 i_1134 (.A(n_580), .B(n_801), .CI(n_692), .CO(n_587), .S(n_586));
   FA_X1 i_1135 (.A(n_582), .B(n_584), .CI(n_828), .CO(n_589), .S(n_588));
   FA_X1 i_1136 (.A(n_583), .B(n_620), .CI(n_585), .CO(n_627), .S(n_626));
   FA_X1 i_1137 (.A(n_622), .B(n_624), .CI(n_587), .CO(n_629), .S(n_628));
   FA_X1 i_1138 (.A(n_626), .B(n_589), .CI(n_628), .CO(n_1750), .S(n_1749));
   FA_X1 i_1139 (.A(n_167), .B(n_461), .CI(n_168), .CO(n_611), .S(n_610));
   FA_X1 i_1140 (.A(n_611), .B(n_648), .CI(n_646), .CO(n_1751), .S(n_656));
   FA_X1 i_1141 (.A(n_771), .B(n_504), .CI(n_169), .CO(n_577), .S(n_576));
   FA_X1 i_1142 (.A(n_535), .B(n_531), .CI(n_527), .CO(n_615), .S(n_614));
   FA_X1 i_1143 (.A(n_547), .B(n_543), .CI(n_539), .CO(n_613), .S(n_612));
   FA_X1 i_1144 (.A(n_577), .B(n_614), .CI(n_612), .CO(n_623), .S(n_622));
   FA_X1 i_1145 (.A(n_549), .B(n_517), .CI(n_513), .CO(n_619), .S(n_618));
   FA_X1 i_1146 (.A(n_523), .B(n_505), .CI(n_565), .CO(n_617), .S(n_616));
   FA_X1 i_1147 (.A(n_619), .B(n_617), .CI(n_654), .CO(n_661), .S(n_660));
   FA_X1 i_1148 (.A(n_656), .B(n_623), .CI(n_660), .CO(n_665), .S(n_664));
   FA_X1 i_1149 (.A(n_697), .B(n_507), .CI(n_690), .CO(n_581), .S(n_580));
   FA_X1 i_1150 (.A(n_616), .B(n_581), .CI(n_618), .CO(n_625), .S(n_624));
   FA_X1 i_1151 (.A(n_509), .B(n_610), .CI(n_521), .CO(n_621), .S(n_620));
   FA_X1 i_1152 (.A(n_615), .B(n_613), .CI(n_650), .CO(n_1752), .S(n_658));
   FA_X1 i_1153 (.A(n_652), .B(n_621), .CI(n_658), .CO(n_663), .S(n_662));
   FA_X1 i_1154 (.A(n_515), .B(n_511), .CI(n_800), .CO(n_583), .S(n_582));
   FA_X1 i_1155 (.A(n_519), .B(n_576), .CI(n_724), .CO(n_585), .S(n_584));
   FA_X1 i_1156 (.A(n_664), .B(n_629), .CI(n_666), .CO(n_1754), .S(n_1753));
   FA_X1 i_1157 (.A(n_1229), .B(n_1252), .CI(n_1275), .CO(n_1755), .S(n_886));
   FA_X1 i_1158 (.A(n_857), .B(n_865), .CI(n_886), .CO(n_1756), .S(n_890));
   FA_X1 i_1159 (.A(n_890), .B(n_873), .CI(n_871), .CO(n_1757), .S(n_896));
   FA_X1 i_1160 (.A(n_1160), .B(n_1183), .CI(n_1206), .CO(n_1758), .S(n_884));
   FA_X1 i_1161 (.A(n_1091), .B(n_1114), .CI(n_1137), .CO(n_1759), .S(n_882));
   FA_X1 i_1162 (.A(n_1022), .B(n_1045), .CI(n_1068), .CO(n_1760), .S(n_880));
   FA_X1 i_1163 (.A(n_884), .B(n_882), .CI(n_880), .CO(n_1761), .S(n_892));
   FA_X1 i_1164 (.A(n_863), .B(n_861), .CI(n_859), .CO(n_1762), .S(n_888));
   FA_X1 i_1165 (.A(n_867), .B(n_888), .CI(n_869), .CO(n_1769), .S(n_894));
   FA_X1 i_1166 (.A(n_892), .B(n_894), .CI(n_875), .CO(n_1770), .S(n_898));
   FA_X1 i_1167 (.A(n_896), .B(n_877), .CI(n_898), .CO(n_1772), .S(n_1771));
   NOR2_X1 i_1168 (.A1(n_1723), .A2(n_1687), .ZN(n_1068));
   NOR2_X1 i_1169 (.A1(n_1686), .A2(n_1724), .ZN(n_1045));
   NOR2_X1 i_1170 (.A1(n_1685), .A2(n_1725), .ZN(n_1022));
   NOR2_X1 i_1171 (.A1(n_1720), .A2(n_1690), .ZN(n_1137));
   NOR2_X1 i_1172 (.A1(n_1721), .A2(n_1689), .ZN(n_1114));
   NOR2_X1 i_1173 (.A1(n_1722), .A2(n_1688), .ZN(n_1091));
   NOR2_X1 i_1174 (.A1(n_1716), .A2(n_1697), .ZN(n_1206));
   NOR2_X1 i_1175 (.A1(n_1718), .A2(n_1696), .ZN(n_1183));
   NOR2_X1 i_1176 (.A1(n_1719), .A2(n_1691), .ZN(n_1160));
   NOR2_X1 i_1177 (.A1(n_1713), .A2(n_1700), .ZN(n_1275));
   NOR2_X1 i_1178 (.A1(n_1699), .A2(n_1714), .ZN(n_1252));
   NOR2_X1 i_1179 (.A1(n_1698), .A2(n_1715), .ZN(n_1229));
   NOR2_X1 i_1180 (.A1(n_1712), .A2(n_1700), .ZN(n_1299));
   NOR2_X1 i_1181 (.A1(n_1716), .A2(n_1696), .ZN(n_1207));
   NOR2_X1 i_1182 (.A1(n_1718), .A2(n_1691), .ZN(n_1184));
   NOR2_X1 i_1183 (.A1(n_1719), .A2(n_1690), .ZN(n_1161));
   NOR2_X1 i_1184 (.A1(n_1699), .A2(n_1713), .ZN(n_1276));
   NOR2_X1 i_1185 (.A1(n_1698), .A2(n_1714), .ZN(n_1253));
   NOR2_X1 i_1186 (.A1(n_1697), .A2(n_1715), .ZN(n_1230));
   NOR2_X1 i_1187 (.A1(n_1686), .A2(n_1723), .ZN(n_1069));
   NOR2_X1 i_1188 (.A1(n_1685), .A2(n_1724), .ZN(n_1046));
   NOR2_X1 i_1189 (.A1(n_1684), .A2(n_1725), .ZN(n_1023));
   NOR2_X1 i_1190 (.A1(n_1720), .A2(n_1689), .ZN(n_1138));
   NOR2_X1 i_1191 (.A1(n_1721), .A2(n_1688), .ZN(n_1115));
   NOR2_X1 i_1192 (.A1(n_1722), .A2(n_1687), .ZN(n_1092));
   NOR2_X1 i_1193 (.A1(n_1700), .A2(n_1706), .ZN(n_1443));
   NOR2_X1 i_1194 (.A1(n_1711), .A2(n_1700), .ZN(n_1323));
   NOR2_X1 i_1195 (.A1(n_1712), .A2(n_1699), .ZN(n_1300));
   NOR2_X1 i_1196 (.A1(n_1710), .A2(n_1700), .ZN(n_1347));
   NOR2_X1 i_1197 (.A1(n_1711), .A2(n_1699), .ZN(n_1324));
   NOR2_X1 i_1198 (.A1(n_1712), .A2(n_1698), .ZN(n_1301));
   NOR2_X1 i_1199 (.A1(n_1684), .A2(n_1723), .ZN(n_1071));
   NOR2_X1 i_1200 (.A1(n_1724), .A2(n_1683), .ZN(n_1048));
   NOR2_X1 i_1201 (.A1(n_1725), .A2(n_1682), .ZN(n_1025));
   NOR2_X1 i_1202 (.A1(n_1723), .A2(n_1679), .ZN(n_1075));
   NOR2_X1 i_1203 (.A1(n_1724), .A2(n_1678), .ZN(n_1052));
   NOR2_X1 i_1204 (.A1(n_1725), .A2(n_1676), .ZN(n_1029));
   NOR2_X1 i_1205 (.A1(n_1720), .A2(n_1683), .ZN(n_1144));
   NOR2_X1 i_1206 (.A1(n_1721), .A2(n_1682), .ZN(n_1121));
   NOR2_X1 i_1207 (.A1(n_1722), .A2(n_1681), .ZN(n_1098));
   NOR2_X1 i_1208 (.A1(n_1686), .A2(n_1716), .ZN(n_1213));
   NOR2_X1 i_1209 (.A1(n_1685), .A2(n_1718), .ZN(n_1190));
   NOR2_X1 i_1210 (.A1(n_1684), .A2(n_1719), .ZN(n_1167));
   NOR2_X1 i_1211 (.A1(n_1681), .A2(n_1723), .ZN(n_1074));
   NOR2_X1 i_1212 (.A1(n_1724), .A2(n_1679), .ZN(n_1051));
   NOR2_X1 i_1213 (.A1(n_1725), .A2(n_1678), .ZN(n_1028));
   NOR2_X1 i_1214 (.A1(n_1684), .A2(n_1720), .ZN(n_1143));
   NOR2_X1 i_1215 (.A1(n_1721), .A2(n_1683), .ZN(n_1120));
   NOR2_X1 i_1216 (.A1(n_1722), .A2(n_1682), .ZN(n_1097));
   NOR2_X1 i_1217 (.A1(n_1713), .A2(n_1689), .ZN(n_1282));
   NOR2_X1 i_1218 (.A1(n_1688), .A2(n_1714), .ZN(n_1259));
   NOR2_X1 i_1219 (.A1(n_1687), .A2(n_1715), .ZN(n_1236));
   NOR2_X1 i_1220 (.A1(n_1710), .A2(n_1696), .ZN(n_1351));
   NOR2_X1 i_1221 (.A1(n_1711), .A2(n_1691), .ZN(n_1328));
   NOR2_X1 i_1222 (.A1(n_1712), .A2(n_1690), .ZN(n_1305));
   NOR2_X1 i_1223 (.A1(n_1699), .A2(n_1707), .ZN(n_1420));
   NOR2_X1 i_1224 (.A1(n_1698), .A2(n_1708), .ZN(n_1397));
   NOR2_X1 i_1225 (.A1(n_1697), .A2(n_1709), .ZN(n_1374));
   NOR2_X1 i_1226 (.A1(n_1691), .A2(n_1713), .ZN(n_1280));
   NOR2_X1 i_1227 (.A1(n_1690), .A2(n_1714), .ZN(n_1257));
   NOR2_X1 i_1228 (.A1(n_1715), .A2(n_1689), .ZN(n_1234));
   NOR2_X1 i_1229 (.A1(n_1698), .A2(n_1710), .ZN(n_1349));
   NOR2_X1 i_1230 (.A1(n_1697), .A2(n_1711), .ZN(n_1326));
   NOR2_X1 i_1231 (.A1(n_1712), .A2(n_1696), .ZN(n_1303));
   NOR2_X1 i_1232 (.A1(n_1709), .A2(n_1700), .ZN(n_1371));
   NOR2_X1 i_1233 (.A1(n_1700), .A2(n_1707), .ZN(n_1419));
   NOR2_X1 i_1234 (.A1(n_1699), .A2(n_1708), .ZN(n_1396));
   NOR2_X1 i_1235 (.A1(n_1698), .A2(n_1709), .ZN(n_1373));
   NOR2_X1 i_1236 (.A1(n_1708), .A2(n_1700), .ZN(n_1395));
   NOR2_X1 i_1237 (.A1(n_1699), .A2(n_1709), .ZN(n_1372));
   NOR2_X1 i_1238 (.A1(n_1687), .A2(n_1716), .ZN(n_1212));
   NOR2_X1 i_1239 (.A1(n_1686), .A2(n_1718), .ZN(n_1189));
   NOR2_X1 i_1240 (.A1(n_1685), .A2(n_1719), .ZN(n_1166));
   NOR2_X1 i_1241 (.A1(n_1690), .A2(n_1713), .ZN(n_1281));
   NOR2_X1 i_1242 (.A1(n_1714), .A2(n_1689), .ZN(n_1258));
   NOR2_X1 i_1243 (.A1(n_1688), .A2(n_1715), .ZN(n_1235));
   NOR2_X1 i_1244 (.A1(n_1697), .A2(n_1710), .ZN(n_1350));
   NOR2_X1 i_1245 (.A1(n_1711), .A2(n_1696), .ZN(n_1327));
   NOR2_X1 i_1246 (.A1(n_1712), .A2(n_1691), .ZN(n_1304));
   NOR2_X1 i_1247 (.A1(n_1720), .A2(n_1687), .ZN(n_1140));
   NOR2_X1 i_1248 (.A1(n_1721), .A2(n_1686), .ZN(n_1117));
   NOR2_X1 i_1249 (.A1(n_1722), .A2(n_1685), .ZN(n_1094));
   NOR2_X1 i_1250 (.A1(n_1716), .A2(n_1690), .ZN(n_1209));
   NOR2_X1 i_1251 (.A1(n_1718), .A2(n_1689), .ZN(n_1186));
   NOR2_X1 i_1252 (.A1(n_1719), .A2(n_1688), .ZN(n_1163));
   NOR2_X1 i_1253 (.A1(n_1697), .A2(n_1713), .ZN(n_1278));
   NOR2_X1 i_1254 (.A1(n_1714), .A2(n_1696), .ZN(n_1255));
   NOR2_X1 i_1255 (.A1(n_1715), .A2(n_1691), .ZN(n_1232));
   NOR2_X1 i_1256 (.A1(n_1685), .A2(n_1723), .ZN(n_1070));
   NOR2_X1 i_1257 (.A1(n_1684), .A2(n_1724), .ZN(n_1047));
   NOR2_X1 i_1258 (.A1(n_1725), .A2(n_1683), .ZN(n_1024));
   NOR2_X1 i_1259 (.A1(n_1720), .A2(n_1688), .ZN(n_1139));
   NOR2_X1 i_1260 (.A1(n_1721), .A2(n_1687), .ZN(n_1116));
   NOR2_X1 i_1261 (.A1(n_1722), .A2(n_1686), .ZN(n_1093));
   NOR2_X1 i_1262 (.A1(n_1716), .A2(n_1691), .ZN(n_1208));
   NOR2_X1 i_1263 (.A1(n_1718), .A2(n_1690), .ZN(n_1185));
   NOR2_X1 i_1264 (.A1(n_1719), .A2(n_1689), .ZN(n_1162));
   NOR2_X1 i_1265 (.A1(n_1698), .A2(n_1713), .ZN(n_1277));
   NOR2_X1 i_1266 (.A1(n_1697), .A2(n_1714), .ZN(n_1254));
   NOR2_X1 i_1267 (.A1(n_1715), .A2(n_1696), .ZN(n_1231));
   NOR2_X1 i_1268 (.A1(n_1716), .A2(n_1689), .ZN(n_1210));
   NOR2_X1 i_1269 (.A1(n_1718), .A2(n_1688), .ZN(n_1187));
   NOR2_X1 i_1270 (.A1(n_1719), .A2(n_1687), .ZN(n_1164));
   NOR2_X1 i_1271 (.A1(n_1713), .A2(n_1696), .ZN(n_1279));
   NOR2_X1 i_1272 (.A1(n_1714), .A2(n_1691), .ZN(n_1256));
   NOR2_X1 i_1273 (.A1(n_1715), .A2(n_1690), .ZN(n_1233));
   NOR2_X1 i_1274 (.A1(n_1710), .A2(n_1699), .ZN(n_1348));
   NOR2_X1 i_1275 (.A1(n_1711), .A2(n_1698), .ZN(n_1325));
   NOR2_X1 i_1276 (.A1(n_1712), .A2(n_1697), .ZN(n_1302));
   NOR2_X1 i_1277 (.A1(n_1682), .A2(n_1723), .ZN(n_1073));
   NOR2_X1 i_1278 (.A1(n_1681), .A2(n_1724), .ZN(n_1050));
   NOR2_X1 i_1279 (.A1(n_1725), .A2(n_1679), .ZN(n_1027));
   NOR2_X1 i_1280 (.A1(n_1685), .A2(n_1720), .ZN(n_1142));
   NOR2_X1 i_1281 (.A1(n_1684), .A2(n_1721), .ZN(n_1119));
   NOR2_X1 i_1282 (.A1(n_1722), .A2(n_1683), .ZN(n_1096));
   NOR2_X1 i_1283 (.A1(n_1716), .A2(n_1688), .ZN(n_1211));
   NOR2_X1 i_1284 (.A1(n_1718), .A2(n_1687), .ZN(n_1188));
   NOR2_X1 i_1285 (.A1(n_1686), .A2(n_1719), .ZN(n_1165));
   NOR2_X1 i_1286 (.A1(n_1723), .A2(n_1683), .ZN(n_1072));
   NOR2_X1 i_1287 (.A1(n_1724), .A2(n_1682), .ZN(n_1049));
   NOR2_X1 i_1288 (.A1(n_1725), .A2(n_1681), .ZN(n_1026));
   NOR2_X1 i_1289 (.A1(n_1720), .A2(n_1686), .ZN(n_1141));
   NOR2_X1 i_1290 (.A1(n_1721), .A2(n_1685), .ZN(n_1118));
   NOR2_X1 i_1291 (.A1(n_1722), .A2(n_1684), .ZN(n_1095));
   XNOR2_X1 i_1292 (.A(n_1778), .B(n_1774), .ZN(mult_res[35]));
   OAI21_X1 i_1293 (.A(n_1776), .B1(n_1735), .B2(n_1771), .ZN(n_1774));
   INV_X1 i_1294 (.A(n_1776), .ZN(n_1775));
   NAND2_X1 i_1295 (.A1(n_1735), .A2(n_1771), .ZN(n_1776));
   NOR2_X1 i_1296 (.A1(n_1735), .A2(n_1771), .ZN(n_1777));
   AOI21_X1 i_1297 (.A(n_1815), .B1(n_1814), .B2(n_1779), .ZN(n_1778));
   INV_X1 i_1298 (.A(n_1780), .ZN(n_1779));
   AOI21_X1 i_1299 (.A(n_1813), .B1(n_1782), .B2(n_1781), .ZN(n_1780));
   NAND2_X1 i_1300 (.A1(n_1732), .A2(n_1740), .ZN(n_1781));
   NOR2_X1 i_1301 (.A1(n_1784), .A2(n_1783), .ZN(n_1782));
   AOI211_X1 i_1302 (.A(n_1803), .B(n_1788), .C1(n_1329), .C2(n_895), .ZN(n_1783));
   OAI221_X1 i_1303 (.A(n_1785), .B1(n_1792), .B2(n_1789), .C1(n_1797), .C2(
      n_1788), .ZN(n_1784));
   INV_X1 i_1304 (.A(n_1786), .ZN(n_1785));
   OAI221_X1 i_1305 (.A(n_1787), .B1(n_1821), .B2(n_1820), .C1(n_1806), .C2(
      n_1791), .ZN(n_1786));
   OAI21_X1 i_1306 (.A(n_1790), .B1(n_1808), .B2(n_1807), .ZN(n_1787));
   OR2_X1 i_1307 (.A1(n_1800), .A2(n_1789), .ZN(n_1788));
   OAI21_X1 i_1308 (.A(n_1790), .B1(n_1745), .B2(n_1746), .ZN(n_1789));
   NOR2_X1 i_1309 (.A1(n_1810), .A2(n_1791), .ZN(n_1790));
   NOR2_X1 i_1310 (.A1(n_1739), .A2(n_1742), .ZN(n_1791));
   AOI222_X1 i_1311 (.A1(n_1744), .A2(n_1754), .B1(n_1819), .B2(n_1794), 
      .C1(n_1801), .C2(n_1793), .ZN(n_1792));
   NAND2_X1 i_1312 (.A1(n_1796), .A2(n_1795), .ZN(n_1793));
   AND2_X1 i_1313 (.A1(n_1750), .A2(n_1753), .ZN(n_1794));
   NAND2_X1 i_1314 (.A1(n_1748), .A2(n_1749), .ZN(n_1795));
   NAND2_X1 i_1315 (.A1(n_1747), .A2(n_855), .ZN(n_1796));
   AOI21_X1 i_1316 (.A(n_1798), .B1(n_684), .B2(n_854), .ZN(n_1797));
   OAI21_X1 i_1317 (.A(n_1799), .B1(n_1585), .B2(n_1584), .ZN(n_1798));
   OAI21_X1 i_1318 (.A(n_1804), .B1(n_1816), .B2(n_1490), .ZN(n_1799));
   OAI21_X1 i_1319 (.A(n_1801), .B1(n_1747), .B2(n_855), .ZN(n_1800));
   NOR3_X1 i_1320 (.A1(n_670), .A2(n_669), .A3(n_668), .ZN(n_1801));
   NOR2_X1 i_1321 (.A1(n_1747), .A2(n_855), .ZN(n_1802));
   NAND2_X1 i_1322 (.A1(n_1513), .A2(n_1804), .ZN(n_1803));
   NOR3_X1 i_1323 (.A1(n_1585), .A2(n_1805), .A3(n_1569), .ZN(n_1804));
   NOR2_X1 i_1324 (.A1(n_878), .A2(n_682), .ZN(n_1805));
   NAND2_X1 i_1325 (.A1(n_1741), .A2(n_1743), .ZN(n_1806));
   AND2_X1 i_1326 (.A1(n_739), .A2(n_770), .ZN(n_1807));
   INV_X1 i_1327 (.A(n_1809), .ZN(n_1808));
   NAND2_X1 i_1328 (.A1(n_1745), .A2(n_1746), .ZN(n_1809));
   OAI21_X1 i_1329 (.A(n_1811), .B1(n_1741), .B2(n_1743), .ZN(n_1810));
   INV_X1 i_1330 (.A(n_1812), .ZN(n_1811));
   NOR2_X1 i_1331 (.A1(n_739), .A2(n_770), .ZN(n_1812));
   NOR2_X1 i_1332 (.A1(n_1732), .A2(n_1740), .ZN(n_1813));
   NAND2_X1 i_1333 (.A1(n_1733), .A2(n_1734), .ZN(n_1814));
   NOR2_X1 i_1334 (.A1(n_1733), .A2(n_1734), .ZN(n_1815));
   INV_X1 i_1335 (.A(n_1536), .ZN(n_1816));
   INV_X1 i_1336 (.A(n_669), .ZN(n_1817));
   INV_X1 i_1337 (.A(n_668), .ZN(n_1818));
   INV_X1 i_1338 (.A(n_670), .ZN(n_1819));
   INV_X1 i_1339 (.A(n_1742), .ZN(n_1820));
   INV_X1 i_1340 (.A(n_1739), .ZN(n_1821));
endmodule

module floating(i_a, i_b, i_clk, o_res);
   input [31:0]i_a;
   input [31:0]i_b;
   input i_clk;
   output [31:0]o_res;

   wire enable;
   wire [2:0]outB;
   wire [2:0]outA;
   wire [31:0]special_res;
   wire [4:0]shamt;
   wire [47:0]mult_res;
   wire Sb;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire b;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire Sa;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire [8:0]E_sum;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_13;
   wire n_0_0_7;
   wire n_0_0_14;
   wire n_0_0_8;
   wire n_0_0_15;
   wire n_0_0_9;
   wire n_0_0_16;
   wire n_0_0_10;
   wire n_0_0_17;
   wire n_0_0_11;
   wire n_0_0_18;
   wire n_0_0_28;
   wire n_0_0_19;
   wire [7:0]Eb;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire [31:0]res;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_205;
   wire n_0_0_208;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_264;
   wire [23:0]Na;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire [23:0]Nb;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_297;
   wire n_0_0_300;
   wire n_0_0_316;
   wire n_0_0_319;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_80;
   wire n_0_0_354;
   wire n_0_84;
   wire n_0_0_356;
   wire n_0_76;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_78;
   wire n_0_0_365;
   wire n_0_0_367;
   wire n_0_82;
   wire n_0_0_368;
   wire n_0_74;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_77;
   wire n_0_0_376;
   wire n_0_0_378;
   wire n_0_81;
   wire n_0_0_379;
   wire n_0_73;
   wire n_0_0_380;
   wire n_0_0_382;
   wire n_0_79;
   wire n_0_0_383;
   wire n_0_0_386;
   wire n_0_0_388;
   wire n_0_83;
   wire n_0_0_389;
   wire n_0_75;
   wire n_0_0_391;
   wire n_0_0_12;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_148;
   wire n_0_0_183;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_231;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_265;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_64;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_62;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_317;
   wire n_0_63;
   wire n_0_0_318;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_325;
   wire n_0_0_328;
   wire n_0_0_331;
   wire n_0_61;
   wire n_0_0_334;
   wire n_0_0_353;
   wire n_0_0_355;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_361;
   wire n_0_0_364;
   wire n_0_0_366;
   wire n_0_0_369;
   wire n_0_0_375;
   wire n_0_0_377;
   wire n_0_0_381;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_69;
   wire n_0_0_387;
   wire n_0_70;
   wire n_0_0_390;
   wire n_0_66;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_65;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_71;
   wire n_0_0_402;
   wire n_0_72;
   wire n_0_0_403;
   wire n_0_68;
   wire n_0_0_404;
   wire n_0_67;

   n_case ncase (.A({Sa, n_0_30, n_0_31, n_0_32, n_0_33, n_0_34, n_0_35, n_0_36, 
      n_0_37, n_0_38, n_0_39, n_0_40, n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, 
      n_0_46, n_0_47, n_0_48, n_0_49, n_0_50, n_0_51, n_0_52, n_0_53, n_0_54, 
      n_0_55, n_0_56, n_0_57, n_0_58, n_0_59, n_0_60}), .B({Sb, n_0_0, n_0_1, 
      n_0_2, n_0_3, n_0_4, n_0_5, n_0_6, b, n_0_7, n_0_8, n_0_9, n_0_10, n_0_11, 
      n_0_12, n_0_13, n_0_14, n_0_15, n_0_16, n_0_17, n_0_18, n_0_19, n_0_20, 
      n_0_21, n_0_22, n_0_23, n_0_24, n_0_25, n_0_26, n_0_27, n_0_28, n_0_29}), 
      .S({special_res[31], special_res[23], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6, special_res[0], uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, 
      uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, 
      uc_25, uc_26, uc_27, uc_28}), .outA(outA), .outB(outB), .enable(enable));
   zero_counter zcn (.M({n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
      n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61}), .Zcount(
      shamt));
   datapath__0_29 i_0_8 (.Nb(Nb), .Na(Na), .mult_res({mult_res[47], mult_res[46], 
      mult_res[45], mult_res[44], mult_res[43], mult_res[42], mult_res[41], 
      mult_res[40], mult_res[39], mult_res[38], mult_res[37], mult_res[36], 
      mult_res[35], mult_res[34], mult_res[33], mult_res[32], mult_res[31], 
      mult_res[30], mult_res[29], mult_res[28], mult_res[27], mult_res[26], 
      mult_res[25], mult_res[24], mult_res[23], uc_29, uc_30, uc_31, uc_32, 
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51}));
   DFF_X1 \o_res_reg[31]  (.D(res[31]), .CK(i_clk), .Q(o_res[31]), .QN());
   DFF_X1 \o_res_reg[30]  (.D(res[30]), .CK(i_clk), .Q(o_res[30]), .QN());
   DFF_X1 \o_res_reg[29]  (.D(res[29]), .CK(i_clk), .Q(o_res[29]), .QN());
   DFF_X1 \o_res_reg[28]  (.D(res[28]), .CK(i_clk), .Q(o_res[28]), .QN());
   DFF_X1 \o_res_reg[27]  (.D(res[27]), .CK(i_clk), .Q(o_res[27]), .QN());
   DFF_X1 \o_res_reg[26]  (.D(res[26]), .CK(i_clk), .Q(o_res[26]), .QN());
   DFF_X1 \o_res_reg[25]  (.D(res[25]), .CK(i_clk), .Q(o_res[25]), .QN());
   DFF_X1 \o_res_reg[24]  (.D(res[24]), .CK(i_clk), .Q(o_res[24]), .QN());
   DFF_X1 \o_res_reg[23]  (.D(res[23]), .CK(i_clk), .Q(o_res[23]), .QN());
   DFF_X1 \o_res_reg[22]  (.D(res[22]), .CK(i_clk), .Q(o_res[22]), .QN());
   DFF_X1 \o_res_reg[21]  (.D(res[21]), .CK(i_clk), .Q(o_res[21]), .QN());
   DFF_X1 \o_res_reg[20]  (.D(res[20]), .CK(i_clk), .Q(o_res[20]), .QN());
   DFF_X1 \o_res_reg[19]  (.D(res[19]), .CK(i_clk), .Q(o_res[19]), .QN());
   DFF_X1 \o_res_reg[18]  (.D(res[18]), .CK(i_clk), .Q(o_res[18]), .QN());
   DFF_X1 \o_res_reg[17]  (.D(res[17]), .CK(i_clk), .Q(o_res[17]), .QN());
   DFF_X1 \o_res_reg[16]  (.D(res[16]), .CK(i_clk), .Q(o_res[16]), .QN());
   DFF_X1 \o_res_reg[15]  (.D(res[15]), .CK(i_clk), .Q(o_res[15]), .QN());
   DFF_X1 \o_res_reg[14]  (.D(res[14]), .CK(i_clk), .Q(o_res[14]), .QN());
   DFF_X1 \o_res_reg[13]  (.D(res[13]), .CK(i_clk), .Q(o_res[13]), .QN());
   DFF_X1 \o_res_reg[12]  (.D(res[12]), .CK(i_clk), .Q(o_res[12]), .QN());
   DFF_X1 \o_res_reg[11]  (.D(res[11]), .CK(i_clk), .Q(o_res[11]), .QN());
   DFF_X1 \o_res_reg[10]  (.D(res[10]), .CK(i_clk), .Q(o_res[10]), .QN());
   DFF_X1 \o_res_reg[9]  (.D(res[9]), .CK(i_clk), .Q(o_res[9]), .QN());
   DFF_X1 \o_res_reg[8]  (.D(res[8]), .CK(i_clk), .Q(o_res[8]), .QN());
   DFF_X1 \o_res_reg[7]  (.D(res[7]), .CK(i_clk), .Q(o_res[7]), .QN());
   DFF_X1 \o_res_reg[6]  (.D(res[6]), .CK(i_clk), .Q(o_res[6]), .QN());
   DFF_X1 \o_res_reg[5]  (.D(res[5]), .CK(i_clk), .Q(o_res[5]), .QN());
   DFF_X1 \o_res_reg[4]  (.D(res[4]), .CK(i_clk), .Q(o_res[4]), .QN());
   DFF_X1 \o_res_reg[3]  (.D(res[3]), .CK(i_clk), .Q(o_res[3]), .QN());
   DFF_X1 \o_res_reg[2]  (.D(res[2]), .CK(i_clk), .Q(o_res[2]), .QN());
   DFF_X1 \o_res_reg[1]  (.D(res[1]), .CK(i_clk), .Q(o_res[1]), .QN());
   DFF_X1 \o_res_reg[0]  (.D(res[0]), .CK(i_clk), .Q(o_res[0]), .QN());
   DFF_X1 \b_reg[31]  (.D(i_b[31]), .CK(i_clk), .Q(Sb), .QN());
   DFF_X1 \b_reg[30]  (.D(i_b[30]), .CK(i_clk), .Q(n_0_0), .QN());
   DFF_X1 \b_reg[29]  (.D(i_b[29]), .CK(i_clk), .Q(n_0_1), .QN());
   DFF_X1 \b_reg[28]  (.D(i_b[28]), .CK(i_clk), .Q(n_0_2), .QN());
   DFF_X1 \b_reg[27]  (.D(i_b[27]), .CK(i_clk), .Q(n_0_3), .QN());
   DFF_X1 \b_reg[26]  (.D(i_b[26]), .CK(i_clk), .Q(n_0_4), .QN());
   DFF_X1 \b_reg[25]  (.D(i_b[25]), .CK(i_clk), .Q(n_0_5), .QN());
   DFF_X1 \b_reg[24]  (.D(i_b[24]), .CK(i_clk), .Q(n_0_6), .QN());
   DFF_X1 \b_reg[23]  (.D(i_b[23]), .CK(i_clk), .Q(b), .QN());
   DFF_X1 \b_reg[22]  (.D(i_b[22]), .CK(i_clk), .Q(n_0_7), .QN());
   DFF_X1 \b_reg[21]  (.D(i_b[21]), .CK(i_clk), .Q(n_0_8), .QN());
   DFF_X1 \b_reg[20]  (.D(i_b[20]), .CK(i_clk), .Q(n_0_9), .QN());
   DFF_X1 \b_reg[19]  (.D(i_b[19]), .CK(i_clk), .Q(n_0_10), .QN());
   DFF_X1 \b_reg[18]  (.D(i_b[18]), .CK(i_clk), .Q(n_0_11), .QN());
   DFF_X1 \b_reg[17]  (.D(i_b[17]), .CK(i_clk), .Q(n_0_12), .QN());
   DFF_X1 \b_reg[16]  (.D(i_b[16]), .CK(i_clk), .Q(n_0_13), .QN());
   DFF_X1 \b_reg[15]  (.D(i_b[15]), .CK(i_clk), .Q(n_0_14), .QN());
   DFF_X1 \b_reg[14]  (.D(i_b[14]), .CK(i_clk), .Q(n_0_15), .QN());
   DFF_X1 \b_reg[13]  (.D(i_b[13]), .CK(i_clk), .Q(n_0_16), .QN());
   DFF_X1 \b_reg[12]  (.D(i_b[12]), .CK(i_clk), .Q(n_0_17), .QN());
   DFF_X1 \b_reg[11]  (.D(i_b[11]), .CK(i_clk), .Q(n_0_18), .QN());
   DFF_X1 \b_reg[10]  (.D(i_b[10]), .CK(i_clk), .Q(n_0_19), .QN());
   DFF_X1 \b_reg[9]  (.D(i_b[9]), .CK(i_clk), .Q(n_0_20), .QN());
   DFF_X1 \b_reg[8]  (.D(i_b[8]), .CK(i_clk), .Q(n_0_21), .QN());
   DFF_X1 \b_reg[7]  (.D(i_b[7]), .CK(i_clk), .Q(n_0_22), .QN());
   DFF_X1 \b_reg[6]  (.D(i_b[6]), .CK(i_clk), .Q(n_0_23), .QN());
   DFF_X1 \b_reg[5]  (.D(i_b[5]), .CK(i_clk), .Q(n_0_24), .QN());
   DFF_X1 \b_reg[4]  (.D(i_b[4]), .CK(i_clk), .Q(n_0_25), .QN());
   DFF_X1 \b_reg[3]  (.D(i_b[3]), .CK(i_clk), .Q(n_0_26), .QN());
   DFF_X1 \b_reg[2]  (.D(i_b[2]), .CK(i_clk), .Q(n_0_27), .QN());
   DFF_X1 \b_reg[1]  (.D(i_b[1]), .CK(i_clk), .Q(n_0_28), .QN());
   DFF_X1 \b_reg[0]  (.D(i_b[0]), .CK(i_clk), .Q(n_0_29), .QN());
   DFF_X1 \a_reg[31]  (.D(i_a[31]), .CK(i_clk), .Q(Sa), .QN());
   DFF_X1 \a_reg[30]  (.D(i_a[30]), .CK(i_clk), .Q(n_0_30), .QN());
   DFF_X1 \a_reg[29]  (.D(i_a[29]), .CK(i_clk), .Q(n_0_31), .QN());
   DFF_X1 \a_reg[28]  (.D(i_a[28]), .CK(i_clk), .Q(n_0_32), .QN());
   DFF_X1 \a_reg[27]  (.D(i_a[27]), .CK(i_clk), .Q(n_0_33), .QN());
   DFF_X1 \a_reg[26]  (.D(i_a[26]), .CK(i_clk), .Q(n_0_34), .QN());
   DFF_X1 \a_reg[25]  (.D(i_a[25]), .CK(i_clk), .Q(n_0_35), .QN());
   DFF_X1 \a_reg[24]  (.D(i_a[24]), .CK(i_clk), .Q(n_0_36), .QN());
   DFF_X1 \a_reg[23]  (.D(i_a[23]), .CK(i_clk), .Q(n_0_37), .QN());
   DFF_X1 \a_reg[22]  (.D(i_a[22]), .CK(i_clk), .Q(n_0_38), .QN());
   DFF_X1 \a_reg[21]  (.D(i_a[21]), .CK(i_clk), .Q(n_0_39), .QN());
   DFF_X1 \a_reg[20]  (.D(i_a[20]), .CK(i_clk), .Q(n_0_40), .QN());
   DFF_X1 \a_reg[19]  (.D(i_a[19]), .CK(i_clk), .Q(n_0_41), .QN());
   DFF_X1 \a_reg[18]  (.D(i_a[18]), .CK(i_clk), .Q(n_0_42), .QN());
   DFF_X1 \a_reg[17]  (.D(i_a[17]), .CK(i_clk), .Q(n_0_43), .QN());
   DFF_X1 \a_reg[16]  (.D(i_a[16]), .CK(i_clk), .Q(n_0_44), .QN());
   DFF_X1 \a_reg[15]  (.D(i_a[15]), .CK(i_clk), .Q(n_0_45), .QN());
   DFF_X1 \a_reg[14]  (.D(i_a[14]), .CK(i_clk), .Q(n_0_46), .QN());
   DFF_X1 \a_reg[13]  (.D(i_a[13]), .CK(i_clk), .Q(n_0_47), .QN());
   DFF_X1 \a_reg[12]  (.D(i_a[12]), .CK(i_clk), .Q(n_0_48), .QN());
   DFF_X1 \a_reg[11]  (.D(i_a[11]), .CK(i_clk), .Q(n_0_49), .QN());
   DFF_X1 \a_reg[10]  (.D(i_a[10]), .CK(i_clk), .Q(n_0_50), .QN());
   DFF_X1 \a_reg[9]  (.D(i_a[9]), .CK(i_clk), .Q(n_0_51), .QN());
   DFF_X1 \a_reg[8]  (.D(i_a[8]), .CK(i_clk), .Q(n_0_52), .QN());
   DFF_X1 \a_reg[7]  (.D(i_a[7]), .CK(i_clk), .Q(n_0_53), .QN());
   DFF_X1 \a_reg[6]  (.D(i_a[6]), .CK(i_clk), .Q(n_0_54), .QN());
   DFF_X1 \a_reg[5]  (.D(i_a[5]), .CK(i_clk), .Q(n_0_55), .QN());
   DFF_X1 \a_reg[4]  (.D(i_a[4]), .CK(i_clk), .Q(n_0_56), .QN());
   DFF_X1 \a_reg[3]  (.D(i_a[3]), .CK(i_clk), .Q(n_0_57), .QN());
   DFF_X1 \a_reg[2]  (.D(i_a[2]), .CK(i_clk), .Q(n_0_58), .QN());
   DFF_X1 \a_reg[1]  (.D(i_a[1]), .CK(i_clk), .Q(n_0_59), .QN());
   DFF_X1 \a_reg[0]  (.D(i_a[0]), .CK(i_clk), .Q(n_0_60), .QN());
   FA_X1 i_0_0_0 (.A(mult_res[47]), .B(n_0_0_34), .CI(Eb[0]), .CO(n_0_0_0), 
      .S(E_sum[0]));
   FA_X1 i_0_0_1 (.A(Eb[1]), .B(n_0_0_32), .CI(n_0_0_0), .CO(n_0_0_1), .S(
      E_sum[1]));
   FA_X1 i_0_0_2 (.A(Eb[2]), .B(n_0_0_30), .CI(n_0_0_1), .CO(n_0_0_2), .S(
      E_sum[2]));
   FA_X1 i_0_0_3 (.A(Eb[3]), .B(n_0_0_69), .CI(n_0_0_2), .CO(n_0_0_3), .S(
      E_sum[3]));
   FA_X1 i_0_0_4 (.A(Eb[4]), .B(n_0_0_25), .CI(n_0_0_3), .CO(n_0_0_4), .S(
      E_sum[4]));
   FA_X1 i_0_0_5 (.A(Eb[5]), .B(n_0_0_23), .CI(n_0_0_4), .CO(n_0_0_5), .S(
      E_sum[5]));
   FA_X1 i_0_0_6 (.A(Eb[6]), .B(n_0_0_21), .CI(n_0_0_5), .CO(n_0_0_6), .S(
      E_sum[6]));
   FA_X1 i_0_0_7 (.A(Eb[7]), .B(n_0_0_19), .CI(n_0_0_6), .CO(E_sum[8]), .S(
      E_sum[7]));
   HA_X1 i_0_0_8 (.A(E_sum[1]), .B(E_sum[0]), .CO(n_0_0_7), .S(n_0_0_13));
   HA_X1 i_0_0_9 (.A(E_sum[2]), .B(n_0_0_7), .CO(n_0_0_8), .S(n_0_0_14));
   HA_X1 i_0_0_10 (.A(E_sum[3]), .B(n_0_0_8), .CO(n_0_0_9), .S(n_0_0_15));
   HA_X1 i_0_0_11 (.A(E_sum[4]), .B(n_0_0_9), .CO(n_0_0_10), .S(n_0_0_16));
   HA_X1 i_0_0_12 (.A(E_sum[5]), .B(n_0_0_10), .CO(n_0_0_11), .S(n_0_0_17));
   HA_X1 i_0_0_13 (.A(E_sum[6]), .B(n_0_0_11), .CO(n_0_0_28), .S(n_0_0_18));
   OAI21_X1 i_0_0_14 (.A(n_0_0_257), .B1(n_0_0_259), .B2(n_0_0_258), .ZN(
      n_0_0_19));
   INV_X1 i_0_0_15 (.A(n_0_0_20), .ZN(Eb[7]));
   AOI22_X1 i_0_0_16 (.A1(n_0_0), .A2(n_0_0_37), .B1(n_0_30), .B2(n_0_0_36), 
      .ZN(n_0_0_20));
   OAI21_X1 i_0_0_17 (.A(n_0_0_260), .B1(n_0_0_262), .B2(n_0_0_261), .ZN(
      n_0_0_21));
   INV_X1 i_0_0_18 (.A(n_0_0_22), .ZN(Eb[6]));
   AOI22_X1 i_0_0_19 (.A1(n_0_1), .A2(n_0_0_37), .B1(n_0_31), .B2(n_0_0_36), 
      .ZN(n_0_0_22));
   OAI21_X1 i_0_0_20 (.A(n_0_0_263), .B1(n_0_0_294), .B2(n_0_0_265), .ZN(
      n_0_0_23));
   INV_X1 i_0_0_21 (.A(n_0_0_24), .ZN(Eb[5]));
   AOI22_X1 i_0_0_22 (.A1(n_0_2), .A2(n_0_0_37), .B1(n_0_32), .B2(n_0_0_36), 
      .ZN(n_0_0_24));
   XOR2_X1 i_0_0_23 (.A(n_0_0_296), .B(n_0_0_26), .Z(n_0_0_25));
   AOI21_X1 i_0_0_24 (.A(n_0_0_299), .B1(shamt[4]), .B2(n_0_0_301), .ZN(n_0_0_26));
   INV_X1 i_0_0_25 (.A(n_0_0_27), .ZN(Eb[4]));
   AOI22_X1 i_0_0_26 (.A1(n_0_3), .A2(n_0_0_37), .B1(n_0_33), .B2(n_0_0_36), 
      .ZN(n_0_0_27));
   INV_X1 i_0_0_27 (.A(n_0_0_29), .ZN(Eb[3]));
   AOI22_X1 i_0_0_28 (.A1(n_0_4), .A2(n_0_0_37), .B1(n_0_34), .B2(n_0_0_36), 
      .ZN(n_0_0_29));
   XNOR2_X1 i_0_0_30 (.A(n_0_0_39), .B(n_0_0_56), .ZN(n_0_0_30));
   INV_X1 i_0_0_31 (.A(n_0_0_31), .ZN(Eb[2]));
   AOI22_X1 i_0_0_32 (.A1(n_0_5), .A2(n_0_0_37), .B1(n_0_35), .B2(n_0_0_36), 
      .ZN(n_0_0_31));
   XNOR2_X1 i_0_0_33 (.A(n_0_0_49), .B(n_0_0_55), .ZN(n_0_0_32));
   INV_X1 i_0_0_34 (.A(n_0_0_33), .ZN(Eb[1]));
   AOI22_X1 i_0_0_35 (.A1(n_0_6), .A2(n_0_0_37), .B1(n_0_36), .B2(n_0_0_36), 
      .ZN(n_0_0_33));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_40), .A2(n_0_84), .ZN(Eb[0]));
   OAI21_X1 i_0_0_37 (.A(n_0_0_49), .B1(shamt[0]), .B2(n_0_0_48), .ZN(n_0_0_34));
   NAND3_X1 i_0_0_36 (.A1(n_0_0_184), .A2(n_0_0_42), .A3(n_0_0_75), .ZN(res[0]));
   NAND2_X1 i_0_0_38 (.A1(mult_res[24]), .A2(n_0_0_185), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_39 (.A1(n_0_0_184), .A2(n_0_0_43), .ZN(res[1]));
   AOI222_X1 i_0_0_40 (.A1(mult_res[25]), .A2(n_0_0_185), .B1(mult_res[24]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_44), .ZN(n_0_0_43));
   AOI22_X1 i_0_0_41 (.A1(E_sum[0]), .A2(n_0_0_52), .B1(n_0_0_302), .B2(n_0_0_94), 
      .ZN(n_0_0_44));
   NAND2_X1 i_0_0_42 (.A1(n_0_0_184), .A2(n_0_0_50), .ZN(res[2]));
   AOI222_X1 i_0_0_43 (.A1(mult_res[26]), .A2(n_0_0_185), .B1(mult_res[25]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_51), .ZN(n_0_0_50));
   AOI22_X1 i_0_0_44 (.A1(E_sum[0]), .A2(n_0_0_59), .B1(n_0_0_302), .B2(n_0_0_52), 
      .ZN(n_0_0_51));
   OAI22_X1 i_0_0_45 (.A1(n_0_0_231), .A2(n_0_0_67), .B1(n_0_0_234), .B2(
      n_0_0_201), .ZN(n_0_0_52));
   NAND2_X1 i_0_0_46 (.A1(n_0_0_184), .A2(n_0_0_57), .ZN(res[3]));
   AOI222_X1 i_0_0_47 (.A1(mult_res[27]), .A2(n_0_0_185), .B1(mult_res[26]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_58), .ZN(n_0_0_57));
   AOI22_X1 i_0_0_48 (.A1(n_0_0_302), .A2(n_0_0_59), .B1(E_sum[0]), .B2(n_0_0_66), 
      .ZN(n_0_0_58));
   OAI22_X1 i_0_0_49 (.A1(n_0_0_231), .A2(n_0_0_74), .B1(n_0_0_234), .B2(
      n_0_0_191), .ZN(n_0_0_59));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_184), .A2(n_0_0_64), .ZN(res[4]));
   AOI222_X1 i_0_0_51 (.A1(mult_res[28]), .A2(n_0_0_185), .B1(mult_res[27]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_65), .ZN(n_0_0_64));
   AOI22_X1 i_0_0_52 (.A1(E_sum[0]), .A2(n_0_0_73), .B1(n_0_0_302), .B2(n_0_0_66), 
      .ZN(n_0_0_65));
   AOI22_X1 i_0_0_53 (.A1(n_0_0_231), .A2(n_0_0_67), .B1(n_0_0_234), .B2(
      n_0_0_83), .ZN(n_0_0_66));
   OAI22_X1 i_0_0_54 (.A1(n_0_0_219), .A2(n_0_0_101), .B1(n_0_0_218), .B2(
      n_0_0_210), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_55 (.A1(n_0_0_184), .A2(n_0_0_71), .ZN(res[5]));
   AOI222_X1 i_0_0_56 (.A1(mult_res[29]), .A2(n_0_0_185), .B1(mult_res[28]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_72), .ZN(n_0_0_71));
   AOI21_X1 i_0_0_57 (.A(n_0_0_78), .B1(n_0_0_302), .B2(n_0_0_73), .ZN(n_0_0_72));
   AOI22_X1 i_0_0_58 (.A1(n_0_0_231), .A2(n_0_0_74), .B1(n_0_0_234), .B2(
      n_0_0_91), .ZN(n_0_0_73));
   OAI22_X1 i_0_0_59 (.A1(n_0_0_218), .A2(n_0_0_198), .B1(n_0_0_219), .B2(
      n_0_0_107), .ZN(n_0_0_74));
   AOI211_X1 i_0_0_60 (.A(n_0_0_82), .B(n_0_0_302), .C1(n_0_0_231), .C2(n_0_0_83), 
      .ZN(n_0_0_78));
   NAND2_X1 i_0_0_61 (.A1(n_0_0_184), .A2(n_0_0_79), .ZN(res[6]));
   AOI222_X1 i_0_0_62 (.A1(mult_res[30]), .A2(n_0_0_185), .B1(mult_res[29]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_80), .ZN(n_0_0_79));
   AOI21_X1 i_0_0_63 (.A(n_0_0_81), .B1(E_sum[0]), .B2(n_0_0_90), .ZN(n_0_0_80));
   AOI211_X1 i_0_0_64 (.A(n_0_0_82), .B(E_sum[0]), .C1(n_0_0_303), .C2(n_0_0_83), 
      .ZN(n_0_0_81));
   AND2_X1 i_0_0_65 (.A1(n_0_0_234), .A2(n_0_0_100), .ZN(n_0_0_82));
   AOI22_X1 i_0_0_66 (.A1(n_0_0_219), .A2(n_0_0_206), .B1(n_0_0_218), .B2(
      n_0_0_114), .ZN(n_0_0_83));
   NAND3_X1 i_0_0_67 (.A1(n_0_0_184), .A2(n_0_0_88), .A3(n_0_0_87), .ZN(res[7]));
   AOI22_X1 i_0_0_68 (.A1(mult_res[31]), .A2(n_0_0_185), .B1(mult_res[30]), 
      .B2(n_0_0_93), .ZN(n_0_0_87));
   OAI21_X1 i_0_0_69 (.A(n_0_0_89), .B1(n_0_0_302), .B2(n_0_0_98), .ZN(n_0_0_88));
   AOI21_X1 i_0_0_70 (.A(n_0_0_190), .B1(n_0_0_302), .B2(n_0_0_90), .ZN(n_0_0_89));
   AOI22_X1 i_0_0_71 (.A1(n_0_0_234), .A2(n_0_0_106), .B1(n_0_0_231), .B2(
      n_0_0_91), .ZN(n_0_0_90));
   OAI22_X1 i_0_0_72 (.A1(n_0_0_218), .A2(n_0_0_195), .B1(n_0_0_219), .B2(
      n_0_0_120), .ZN(n_0_0_91));
   NAND2_X1 i_0_0_73 (.A1(n_0_0_184), .A2(n_0_0_95), .ZN(res[8]));
   AOI222_X1 i_0_0_74 (.A1(mult_res[32]), .A2(n_0_0_185), .B1(mult_res[31]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_96), .ZN(n_0_0_95));
   OAI21_X1 i_0_0_75 (.A(n_0_0_97), .B1(n_0_0_302), .B2(n_0_0_105), .ZN(n_0_0_96));
   NAND2_X1 i_0_0_76 (.A1(n_0_0_302), .A2(n_0_0_98), .ZN(n_0_0_97));
   AOI21_X1 i_0_0_77 (.A(n_0_0_99), .B1(n_0_0_234), .B2(n_0_0_112), .ZN(n_0_0_98));
   NOR2_X1 i_0_0_78 (.A1(n_0_0_234), .A2(n_0_0_100), .ZN(n_0_0_99));
   AOI22_X1 i_0_0_79 (.A1(n_0_0_219), .A2(n_0_0_101), .B1(n_0_0_218), .B2(
      n_0_0_127), .ZN(n_0_0_100));
   AOI22_X1 i_0_0_80 (.A1(mult_res[31]), .A2(n_0_0_208), .B1(mult_res[39]), 
      .B2(n_0_0_213), .ZN(n_0_0_101));
   NAND3_X1 i_0_0_81 (.A1(n_0_0_184), .A2(n_0_0_103), .A3(n_0_0_102), .ZN(res[9]));
   AOI22_X1 i_0_0_82 (.A1(mult_res[33]), .A2(n_0_0_185), .B1(mult_res[32]), 
      .B2(n_0_0_93), .ZN(n_0_0_102));
   OAI21_X1 i_0_0_83 (.A(n_0_0_104), .B1(n_0_0_302), .B2(n_0_0_111), .ZN(
      n_0_0_103));
   AOI21_X1 i_0_0_84 (.A(n_0_0_190), .B1(n_0_0_302), .B2(n_0_0_105), .ZN(
      n_0_0_104));
   AOI22_X1 i_0_0_85 (.A1(n_0_0_231), .A2(n_0_0_106), .B1(n_0_0_234), .B2(
      n_0_0_119), .ZN(n_0_0_105));
   OAI22_X1 i_0_0_86 (.A1(n_0_0_219), .A2(n_0_0_133), .B1(n_0_0_218), .B2(
      n_0_0_107), .ZN(n_0_0_106));
   AOI22_X1 i_0_0_87 (.A1(mult_res[32]), .A2(n_0_0_208), .B1(mult_res[40]), 
      .B2(n_0_0_213), .ZN(n_0_0_107));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_184), .A2(n_0_0_108), .ZN(res[10]));
   AOI222_X1 i_0_0_122 (.A1(mult_res[34]), .A2(n_0_0_185), .B1(mult_res[33]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_109), .ZN(n_0_0_108));
   OAI21_X1 i_0_0_123 (.A(n_0_0_110), .B1(n_0_0_302), .B2(n_0_0_118), .ZN(
      n_0_0_109));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_302), .A2(n_0_0_111), .ZN(n_0_0_110));
   AOI22_X1 i_0_0_88 (.A1(n_0_0_231), .A2(n_0_0_112), .B1(n_0_0_234), .B2(
      n_0_0_125), .ZN(n_0_0_111));
   OAI21_X1 i_0_0_89 (.A(n_0_0_113), .B1(n_0_0_219), .B2(n_0_0_140), .ZN(
      n_0_0_112));
   NAND2_X1 i_0_0_90 (.A1(n_0_0_219), .A2(n_0_0_114), .ZN(n_0_0_113));
   AOI22_X1 i_0_0_91 (.A1(mult_res[33]), .A2(n_0_0_208), .B1(mult_res[41]), 
      .B2(n_0_0_213), .ZN(n_0_0_114));
   NAND3_X1 i_0_0_129 (.A1(n_0_0_184), .A2(n_0_0_116), .A3(n_0_0_115), .ZN(
      res[11]));
   AOI22_X1 i_0_0_130 (.A1(mult_res[35]), .A2(n_0_0_185), .B1(mult_res[34]), 
      .B2(n_0_0_93), .ZN(n_0_0_115));
   OAI21_X1 i_0_0_131 (.A(n_0_0_117), .B1(n_0_0_302), .B2(n_0_0_124), .ZN(
      n_0_0_116));
   AOI21_X1 i_0_0_132 (.A(n_0_0_190), .B1(n_0_0_302), .B2(n_0_0_118), .ZN(
      n_0_0_117));
   AOI22_X1 i_0_0_133 (.A1(n_0_0_231), .A2(n_0_0_119), .B1(n_0_0_234), .B2(
      n_0_0_132), .ZN(n_0_0_118));
   OAI22_X1 i_0_0_92 (.A1(n_0_0_219), .A2(n_0_0_147), .B1(n_0_0_218), .B2(
      n_0_0_120), .ZN(n_0_0_119));
   AOI22_X1 i_0_0_93 (.A1(mult_res[34]), .A2(n_0_0_208), .B1(mult_res[42]), 
      .B2(n_0_0_213), .ZN(n_0_0_120));
   NAND2_X1 i_0_0_136 (.A1(n_0_0_184), .A2(n_0_0_121), .ZN(res[12]));
   AOI222_X1 i_0_0_137 (.A1(mult_res[36]), .A2(n_0_0_185), .B1(mult_res[35]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_122), .ZN(n_0_0_121));
   OAI21_X1 i_0_0_138 (.A(n_0_0_123), .B1(n_0_0_302), .B2(n_0_0_131), .ZN(
      n_0_0_122));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_302), .A2(n_0_0_124), .ZN(n_0_0_123));
   AOI22_X1 i_0_0_140 (.A1(n_0_0_231), .A2(n_0_0_125), .B1(n_0_0_234), .B2(
      n_0_0_139), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_94 (.A1(n_0_0_219), .A2(n_0_0_126), .B1(mult_res[39]), 
      .B2(n_0_0_173), .ZN(n_0_0_125));
   INV_X1 i_0_0_95 (.A(n_0_0_127), .ZN(n_0_0_126));
   AOI22_X1 i_0_0_96 (.A1(mult_res[35]), .A2(n_0_0_208), .B1(mult_res[43]), 
      .B2(n_0_0_213), .ZN(n_0_0_127));
   NAND3_X1 i_0_0_144 (.A1(n_0_0_184), .A2(n_0_0_129), .A3(n_0_0_128), .ZN(
      res[13]));
   AOI22_X1 i_0_0_145 (.A1(mult_res[37]), .A2(n_0_0_185), .B1(mult_res[36]), 
      .B2(n_0_0_93), .ZN(n_0_0_128));
   OAI21_X1 i_0_0_146 (.A(n_0_0_130), .B1(n_0_0_302), .B2(n_0_0_138), .ZN(
      n_0_0_129));
   AOI21_X1 i_0_0_147 (.A(n_0_0_190), .B1(n_0_0_302), .B2(n_0_0_131), .ZN(
      n_0_0_130));
   AOI22_X1 i_0_0_148 (.A1(n_0_0_231), .A2(n_0_0_132), .B1(n_0_0_234), .B2(
      n_0_0_146), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_149 (.A(n_0_0_134), .B1(n_0_0_218), .B2(n_0_0_133), .ZN(
      n_0_0_132));
   AOI22_X1 i_0_0_97 (.A1(mult_res[36]), .A2(n_0_0_208), .B1(mult_res[44]), 
      .B2(n_0_0_213), .ZN(n_0_0_133));
   NAND2_X1 i_0_0_151 (.A1(mult_res[40]), .A2(n_0_0_173), .ZN(n_0_0_134));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_184), .A2(n_0_0_135), .ZN(res[14]));
   AOI221_X1 i_0_0_153 (.A(n_0_0_136), .B1(mult_res[38]), .B2(n_0_0_185), 
      .C1(mult_res[37]), .C2(n_0_0_93), .ZN(n_0_0_135));
   AOI221_X1 i_0_0_154 (.A(n_0_0_190), .B1(E_sum[0]), .B2(n_0_0_145), .C1(
      n_0_0_302), .C2(n_0_0_137), .ZN(n_0_0_136));
   INV_X1 i_0_0_155 (.A(n_0_0_138), .ZN(n_0_0_137));
   AOI22_X1 i_0_0_156 (.A1(n_0_0_234), .A2(n_0_0_154), .B1(n_0_0_231), .B2(
      n_0_0_139), .ZN(n_0_0_138));
   AOI22_X1 i_0_0_157 (.A1(n_0_0_219), .A2(n_0_0_140), .B1(mult_res[41]), 
      .B2(n_0_0_173), .ZN(n_0_0_139));
   INV_X1 i_0_0_98 (.A(n_0_0_141), .ZN(n_0_0_140));
   AOI22_X1 i_0_0_99 (.A1(mult_res[37]), .A2(n_0_0_208), .B1(mult_res[45]), 
      .B2(n_0_0_213), .ZN(n_0_0_141));
   NAND3_X1 i_0_0_160 (.A1(n_0_0_184), .A2(n_0_0_143), .A3(n_0_0_142), .ZN(
      res[15]));
   AOI22_X1 i_0_0_161 (.A1(mult_res[39]), .A2(n_0_0_185), .B1(mult_res[38]), 
      .B2(n_0_0_93), .ZN(n_0_0_142));
   OAI21_X1 i_0_0_162 (.A(n_0_0_144), .B1(n_0_0_302), .B2(n_0_0_153), .ZN(
      n_0_0_143));
   AOI21_X1 i_0_0_163 (.A(n_0_0_190), .B1(n_0_0_302), .B2(n_0_0_145), .ZN(
      n_0_0_144));
   AOI22_X1 i_0_0_100 (.A1(n_0_0_231), .A2(n_0_0_146), .B1(n_0_0_234), .B2(
      n_0_0_158), .ZN(n_0_0_145));
   OAI21_X1 i_0_0_101 (.A(n_0_0_149), .B1(n_0_0_218), .B2(n_0_0_147), .ZN(
      n_0_0_146));
   AOI22_X1 i_0_0_102 (.A1(mult_res[38]), .A2(n_0_0_208), .B1(mult_res[46]), 
      .B2(n_0_0_213), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_103 (.A1(mult_res[42]), .A2(n_0_0_173), .ZN(n_0_0_149));
   NAND3_X1 i_0_0_104 (.A1(n_0_0_184), .A2(n_0_0_151), .A3(n_0_0_150), .ZN(
      res[16]));
   AOI22_X1 i_0_0_105 (.A1(mult_res[40]), .A2(n_0_0_185), .B1(mult_res[39]), 
      .B2(n_0_0_93), .ZN(n_0_0_150));
   OAI21_X1 i_0_0_106 (.A(n_0_0_152), .B1(E_sum[0]), .B2(n_0_0_153), .ZN(
      n_0_0_151));
   AOI21_X1 i_0_0_107 (.A(n_0_0_190), .B1(E_sum[0]), .B2(n_0_0_157), .ZN(
      n_0_0_152));
   AOI22_X1 i_0_0_108 (.A1(n_0_0_231), .A2(n_0_0_154), .B1(n_0_0_234), .B2(
      n_0_0_165), .ZN(n_0_0_153));
   AOI22_X1 i_0_0_109 (.A1(mult_res[43]), .A2(n_0_0_173), .B1(mult_res[39]), 
      .B2(n_0_0_205), .ZN(n_0_0_154));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_184), .A2(n_0_0_155), .ZN(res[17]));
   AOI221_X1 i_0_0_176 (.A(n_0_0_156), .B1(mult_res[41]), .B2(n_0_0_185), 
      .C1(mult_res[40]), .C2(n_0_0_93), .ZN(n_0_0_155));
   AOI221_X1 i_0_0_177 (.A(n_0_0_190), .B1(E_sum[0]), .B2(n_0_0_162), .C1(
      n_0_0_302), .C2(n_0_0_157), .ZN(n_0_0_156));
   AOI22_X1 i_0_0_110 (.A1(n_0_0_231), .A2(n_0_0_158), .B1(n_0_0_234), .B2(
      n_0_0_171), .ZN(n_0_0_157));
   INV_X1 i_0_0_111 (.A(n_0_0_159), .ZN(n_0_0_158));
   AOI22_X1 i_0_0_112 (.A1(mult_res[44]), .A2(n_0_0_173), .B1(mult_res[40]), 
      .B2(n_0_0_205), .ZN(n_0_0_159));
   NAND2_X1 i_0_0_181 (.A1(n_0_0_184), .A2(n_0_0_160), .ZN(res[18]));
   AOI221_X1 i_0_0_182 (.A(n_0_0_161), .B1(mult_res[42]), .B2(n_0_0_185), 
      .C1(mult_res[41]), .C2(n_0_0_93), .ZN(n_0_0_160));
   AOI221_X1 i_0_0_183 (.A(n_0_0_190), .B1(E_sum[0]), .B2(n_0_0_169), .C1(
      n_0_0_302), .C2(n_0_0_162), .ZN(n_0_0_161));
   INV_X1 i_0_0_184 (.A(n_0_0_163), .ZN(n_0_0_162));
   OAI21_X1 i_0_0_185 (.A(n_0_0_164), .B1(n_0_0_234), .B2(n_0_0_165), .ZN(
      n_0_0_163));
   NAND3_X1 i_0_0_186 (.A1(mult_res[43]), .A2(n_0_0_205), .A3(n_0_0_234), 
      .ZN(n_0_0_164));
   AOI22_X1 i_0_0_113 (.A1(mult_res[45]), .A2(n_0_0_173), .B1(mult_res[41]), 
      .B2(n_0_0_205), .ZN(n_0_0_165));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_184), .A2(n_0_0_166), .ZN(res[19]));
   AOI222_X1 i_0_0_189 (.A1(mult_res[43]), .A2(n_0_0_185), .B1(mult_res[42]), 
      .B2(n_0_0_93), .C1(n_0_0_235), .C2(n_0_0_167), .ZN(n_0_0_166));
   AOI21_X1 i_0_0_190 (.A(n_0_0_168), .B1(n_0_0_302), .B2(n_0_0_169), .ZN(
      n_0_0_167));
   AOI21_X1 i_0_0_191 (.A(n_0_0_302), .B1(n_0_0_205), .B2(n_0_0_176), .ZN(
      n_0_0_168));
   AOI21_X1 i_0_0_192 (.A(n_0_0_170), .B1(n_0_0_231), .B2(n_0_0_171), .ZN(
      n_0_0_169));
   AND3_X1 i_0_0_193 (.A1(mult_res[44]), .A2(n_0_0_205), .A3(n_0_0_234), 
      .ZN(n_0_0_170));
   INV_X1 i_0_0_114 (.A(n_0_0_172), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_115 (.A1(mult_res[46]), .A2(n_0_0_173), .B1(mult_res[42]), 
      .B2(n_0_0_205), .ZN(n_0_0_172));
   AND2_X1 i_0_0_116 (.A1(n_0_0_208), .A2(n_0_0_218), .ZN(n_0_0_173));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_184), .A2(n_0_0_174), .ZN(res[20]));
   AOI222_X1 i_0_0_198 (.A1(n_0_0_189), .A2(n_0_0_175), .B1(mult_res[44]), 
      .B2(n_0_0_185), .C1(mult_res[43]), .C2(n_0_0_93), .ZN(n_0_0_174));
   OAI22_X1 i_0_0_199 (.A1(E_sum[0]), .A2(n_0_0_177), .B1(n_0_0_302), .B2(
      n_0_0_181), .ZN(n_0_0_175));
   INV_X1 i_0_0_200 (.A(n_0_0_177), .ZN(n_0_0_176));
   OAI22_X1 i_0_0_201 (.A1(mult_res[45]), .A2(n_0_0_231), .B1(mult_res[43]), 
      .B2(n_0_0_234), .ZN(n_0_0_177));
   NAND2_X1 i_0_0_202 (.A1(n_0_0_184), .A2(n_0_0_178), .ZN(res[21]));
   AOI222_X1 i_0_0_203 (.A1(mult_res[44]), .A2(n_0_0_93), .B1(mult_res[45]), 
      .B2(n_0_0_185), .C1(n_0_0_189), .C2(n_0_0_179), .ZN(n_0_0_178));
   AOI21_X1 i_0_0_204 (.A(n_0_0_180), .B1(n_0_0_302), .B2(n_0_0_181), .ZN(
      n_0_0_179));
   AOI21_X1 i_0_0_205 (.A(n_0_0_302), .B1(mult_res[45]), .B2(E_sum[1]), .ZN(
      n_0_0_180));
   AOI22_X1 i_0_0_206 (.A1(mult_res[44]), .A2(n_0_0_231), .B1(mult_res[46]), 
      .B2(n_0_0_234), .ZN(n_0_0_181));
   OAI211_X1 i_0_0_207 (.A(n_0_0_184), .B(n_0_0_182), .C1(n_0_0_234), .C2(
      n_0_0_186), .ZN(res[22]));
   AOI22_X1 i_0_0_208 (.A1(mult_res[46]), .A2(n_0_0_185), .B1(mult_res[45]), 
      .B2(n_0_0_93), .ZN(n_0_0_182));
   NAND2_X1 i_0_0_117 (.A1(special_res[0]), .A2(n_0_0_309), .ZN(n_0_0_184));
   NOR3_X1 i_0_0_118 (.A1(n_0_0_12), .A2(n_0_0_248), .A3(n_0_0_242), .ZN(
      n_0_0_185));
   OAI221_X1 i_0_0_212 (.A(n_0_0_189), .B1(mult_res[46]), .B2(n_0_0_303), 
      .C1(mult_res[45]), .C2(E_sum[0]), .ZN(n_0_0_186));
   AND2_X1 i_0_0_215 (.A1(n_0_0_205), .A2(n_0_0_235), .ZN(n_0_0_189));
   INV_X1 i_0_0_119 (.A(n_0_0_235), .ZN(n_0_0_190));
   NOR3_X1 i_0_0_120 (.A1(n_0_0_217), .A2(n_0_0_214), .A3(n_0_0_218), .ZN(
      n_0_0_205));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_217), .A2(n_0_0_214), .ZN(n_0_0_208));
   INV_X1 i_0_0_126 (.A(n_0_0_220), .ZN(res[23]));
   AOI21_X1 i_0_0_127 (.A(n_0_0_232), .B1(n_0_0_302), .B2(n_0_0_230), .ZN(
      n_0_0_220));
   INV_X1 i_0_0_248 (.A(n_0_0_221), .ZN(res[24]));
   AOI21_X1 i_0_0_249 (.A(n_0_0_232), .B1(n_0_0_13), .B2(n_0_0_230), .ZN(
      n_0_0_221));
   INV_X1 i_0_0_250 (.A(n_0_0_222), .ZN(res[25]));
   AOI21_X1 i_0_0_251 (.A(n_0_0_232), .B1(n_0_0_14), .B2(n_0_0_230), .ZN(
      n_0_0_222));
   INV_X1 i_0_0_252 (.A(n_0_0_223), .ZN(res[26]));
   AOI21_X1 i_0_0_253 (.A(n_0_0_232), .B1(n_0_0_15), .B2(n_0_0_230), .ZN(
      n_0_0_223));
   INV_X1 i_0_0_254 (.A(n_0_0_224), .ZN(res[27]));
   AOI21_X1 i_0_0_255 (.A(n_0_0_232), .B1(n_0_0_16), .B2(n_0_0_230), .ZN(
      n_0_0_224));
   INV_X1 i_0_0_256 (.A(n_0_0_225), .ZN(res[28]));
   AOI21_X1 i_0_0_257 (.A(n_0_0_232), .B1(n_0_0_17), .B2(n_0_0_230), .ZN(
      n_0_0_225));
   INV_X1 i_0_0_258 (.A(n_0_0_226), .ZN(res[29]));
   AOI21_X1 i_0_0_259 (.A(n_0_0_232), .B1(n_0_0_18), .B2(n_0_0_230), .ZN(
      n_0_0_226));
   INV_X1 i_0_0_260 (.A(n_0_0_227), .ZN(res[30]));
   AOI21_X1 i_0_0_261 (.A(n_0_0_232), .B1(n_0_0_230), .B2(n_0_0_228), .ZN(
      n_0_0_227));
   INV_X1 i_0_0_262 (.A(n_0_0_229), .ZN(n_0_0_228));
   AOI21_X1 i_0_0_263 (.A(n_0_0_256), .B1(E_sum[7]), .B2(n_0_0_28), .ZN(
      n_0_0_229));
   NOR2_X1 i_0_0_128 (.A1(n_0_0_309), .A2(n_0_0_247), .ZN(n_0_0_230));
   OAI21_X1 i_0_0_134 (.A(n_0_0_264), .B1(n_0_0_309), .B2(n_0_0_233), .ZN(
      n_0_0_232));
   NAND3_X1 i_0_0_135 (.A1(E_sum[8]), .A2(n_0_0_255), .A3(n_0_0_257), .ZN(
      n_0_0_233));
   NAND2_X1 i_0_0_141 (.A1(special_res[23]), .A2(n_0_0_309), .ZN(n_0_0_264));
   INV_X1 i_0_0_301 (.A(n_0_0_266), .ZN(Na[0]));
   AOI22_X1 i_0_0_302 (.A1(n_0_60), .A2(n_0_0_37), .B1(n_0_29), .B2(n_0_0_36), 
      .ZN(n_0_0_266));
   INV_X1 i_0_0_303 (.A(n_0_0_267), .ZN(Na[1]));
   AOI22_X1 i_0_0_304 (.A1(n_0_59), .A2(n_0_0_37), .B1(n_0_28), .B2(n_0_0_36), 
      .ZN(n_0_0_267));
   INV_X1 i_0_0_305 (.A(n_0_0_268), .ZN(Na[2]));
   AOI22_X1 i_0_0_306 (.A1(n_0_58), .A2(n_0_0_37), .B1(n_0_27), .B2(n_0_0_36), 
      .ZN(n_0_0_268));
   INV_X1 i_0_0_307 (.A(n_0_0_269), .ZN(Na[3]));
   AOI22_X1 i_0_0_308 (.A1(n_0_57), .A2(n_0_0_37), .B1(n_0_26), .B2(n_0_0_36), 
      .ZN(n_0_0_269));
   INV_X1 i_0_0_309 (.A(n_0_0_270), .ZN(Na[4]));
   AOI22_X1 i_0_0_310 (.A1(n_0_56), .A2(n_0_0_37), .B1(n_0_25), .B2(n_0_0_36), 
      .ZN(n_0_0_270));
   INV_X1 i_0_0_311 (.A(n_0_0_271), .ZN(Na[5]));
   AOI22_X1 i_0_0_312 (.A1(n_0_55), .A2(n_0_0_37), .B1(n_0_24), .B2(n_0_0_36), 
      .ZN(n_0_0_271));
   INV_X1 i_0_0_313 (.A(n_0_0_272), .ZN(Na[6]));
   AOI22_X1 i_0_0_314 (.A1(n_0_54), .A2(n_0_0_37), .B1(n_0_23), .B2(n_0_0_36), 
      .ZN(n_0_0_272));
   INV_X1 i_0_0_315 (.A(n_0_0_273), .ZN(Na[7]));
   AOI22_X1 i_0_0_316 (.A1(n_0_53), .A2(n_0_0_37), .B1(n_0_22), .B2(n_0_0_36), 
      .ZN(n_0_0_273));
   INV_X1 i_0_0_317 (.A(n_0_0_274), .ZN(Na[8]));
   AOI22_X1 i_0_0_318 (.A1(n_0_52), .A2(n_0_0_37), .B1(n_0_21), .B2(n_0_0_36), 
      .ZN(n_0_0_274));
   INV_X1 i_0_0_319 (.A(n_0_0_275), .ZN(Na[9]));
   AOI22_X1 i_0_0_320 (.A1(n_0_51), .A2(n_0_0_37), .B1(n_0_20), .B2(n_0_0_36), 
      .ZN(n_0_0_275));
   INV_X1 i_0_0_321 (.A(n_0_0_276), .ZN(Na[10]));
   AOI22_X1 i_0_0_322 (.A1(n_0_50), .A2(n_0_0_37), .B1(n_0_19), .B2(n_0_0_36), 
      .ZN(n_0_0_276));
   INV_X1 i_0_0_323 (.A(n_0_0_277), .ZN(Na[11]));
   AOI22_X1 i_0_0_324 (.A1(n_0_49), .A2(n_0_0_37), .B1(n_0_18), .B2(n_0_0_36), 
      .ZN(n_0_0_277));
   INV_X1 i_0_0_325 (.A(n_0_0_278), .ZN(Na[12]));
   AOI22_X1 i_0_0_326 (.A1(n_0_48), .A2(n_0_0_37), .B1(n_0_17), .B2(n_0_0_36), 
      .ZN(n_0_0_278));
   INV_X1 i_0_0_327 (.A(n_0_0_279), .ZN(Na[13]));
   AOI22_X1 i_0_0_328 (.A1(n_0_47), .A2(n_0_0_37), .B1(n_0_16), .B2(n_0_0_36), 
      .ZN(n_0_0_279));
   INV_X1 i_0_0_329 (.A(n_0_0_280), .ZN(Na[14]));
   AOI22_X1 i_0_0_330 (.A1(n_0_46), .A2(n_0_0_37), .B1(n_0_15), .B2(n_0_0_36), 
      .ZN(n_0_0_280));
   INV_X1 i_0_0_331 (.A(n_0_0_281), .ZN(Na[15]));
   AOI22_X1 i_0_0_332 (.A1(n_0_45), .A2(n_0_0_37), .B1(n_0_14), .B2(n_0_0_36), 
      .ZN(n_0_0_281));
   INV_X1 i_0_0_333 (.A(n_0_0_282), .ZN(Na[16]));
   AOI22_X1 i_0_0_334 (.A1(n_0_44), .A2(n_0_0_37), .B1(n_0_13), .B2(n_0_0_36), 
      .ZN(n_0_0_282));
   INV_X1 i_0_0_335 (.A(n_0_0_283), .ZN(Na[17]));
   AOI22_X1 i_0_0_336 (.A1(n_0_43), .A2(n_0_0_37), .B1(n_0_12), .B2(n_0_0_36), 
      .ZN(n_0_0_283));
   INV_X1 i_0_0_337 (.A(n_0_0_284), .ZN(Na[18]));
   AOI22_X1 i_0_0_338 (.A1(n_0_42), .A2(n_0_0_37), .B1(n_0_11), .B2(n_0_0_36), 
      .ZN(n_0_0_284));
   INV_X1 i_0_0_339 (.A(n_0_0_285), .ZN(Na[19]));
   AOI22_X1 i_0_0_340 (.A1(n_0_41), .A2(n_0_0_37), .B1(n_0_10), .B2(n_0_0_36), 
      .ZN(n_0_0_285));
   INV_X1 i_0_0_341 (.A(n_0_0_286), .ZN(Na[20]));
   AOI22_X1 i_0_0_342 (.A1(n_0_40), .A2(n_0_0_37), .B1(n_0_9), .B2(n_0_0_36), 
      .ZN(n_0_0_286));
   INV_X1 i_0_0_343 (.A(n_0_0_287), .ZN(Na[21]));
   AOI22_X1 i_0_0_344 (.A1(n_0_39), .A2(n_0_0_37), .B1(n_0_8), .B2(n_0_0_36), 
      .ZN(n_0_0_287));
   INV_X1 i_0_0_345 (.A(n_0_0_288), .ZN(Na[22]));
   AOI22_X1 i_0_0_346 (.A1(n_0_38), .A2(n_0_0_37), .B1(n_0_7), .B2(n_0_0_36), 
      .ZN(n_0_0_288));
   NAND2_X1 i_0_0_347 (.A1(n_0_0_36), .A2(n_0_0_45), .ZN(Na[23]));
   AND3_X1 i_0_0_142 (.A1(n_0_0_353), .A2(n_0_0_293), .A3(n_0_61), .ZN(Nb[0]));
   OAI21_X1 i_0_0_143 (.A(n_0_0_289), .B1(n_0_0_334), .B2(n_0_0_290), .ZN(Nb[1]));
   NAND3_X1 i_0_0_150 (.A1(n_0_0_353), .A2(n_0_0_293), .A3(n_0_62), .ZN(
      n_0_0_289));
   OAI22_X1 i_0_0_158 (.A1(shamt[0]), .A2(n_0_0_291), .B1(n_0_0_314), .B2(
      n_0_0_290), .ZN(Nb[2]));
   NAND2_X1 i_0_0_159 (.A1(shamt[0]), .A2(n_0_0_293), .ZN(n_0_0_290));
   AOI22_X1 i_0_0_164 (.A1(n_0_0_353), .A2(n_0_0_292), .B1(shamt[0]), .B2(
      n_0_0_291), .ZN(Nb[3]));
   AOI22_X1 i_0_0_165 (.A1(n_0_63), .A2(n_0_0_293), .B1(n_0_61), .B2(n_0_0_317), 
      .ZN(n_0_0_291));
   OAI22_X1 i_0_0_166 (.A1(n_0_0_353), .A2(n_0_0_292), .B1(shamt[0]), .B2(
      n_0_0_315), .ZN(Nb[4]));
   AOI22_X1 i_0_0_167 (.A1(n_0_62), .A2(n_0_0_317), .B1(n_0_64), .B2(n_0_0_293), 
      .ZN(n_0_0_292));
   NOR2_X1 i_0_0_168 (.A1(shamt[1]), .A2(n_0_0_321), .ZN(n_0_0_293));
   OAI22_X1 i_0_0_169 (.A1(n_0_0_353), .A2(n_0_0_310), .B1(shamt[0]), .B2(
      n_0_0_297), .ZN(Nb[6]));
   OAI22_X1 i_0_0_170 (.A1(n_0_0_353), .A2(n_0_0_297), .B1(shamt[0]), .B2(
      n_0_0_300), .ZN(Nb[7]));
   AOI22_X1 i_0_0_171 (.A1(shamt[1]), .A2(n_0_0_320), .B1(n_0_0_355), .B2(
      n_0_0_375), .ZN(n_0_0_297));
   OAI22_X1 i_0_0_172 (.A1(n_0_0_353), .A2(n_0_0_300), .B1(shamt[0]), .B2(
      n_0_0_369), .ZN(Nb[8]));
   AOI22_X1 i_0_0_173 (.A1(shamt[1]), .A2(n_0_0_312), .B1(n_0_0_355), .B2(
      n_0_0_358), .ZN(n_0_0_300));
   OAI22_X1 i_0_0_174 (.A1(n_0_0_353), .A2(n_0_0_357), .B1(shamt[0]), .B2(
      n_0_0_399), .ZN(Nb[10]));
   OAI22_X1 i_0_0_178 (.A1(n_0_0_353), .A2(n_0_0_396), .B1(shamt[0]), .B2(
      n_0_0_316), .ZN(Nb[12]));
   OAI22_X1 i_0_0_179 (.A1(n_0_0_353), .A2(n_0_0_316), .B1(shamt[0]), .B2(
      n_0_0_319), .ZN(Nb[13]));
   AOI22_X1 i_0_0_180 (.A1(shamt[1]), .A2(n_0_0_400), .B1(n_0_0_355), .B2(
      n_0_0_324), .ZN(n_0_0_316));
   OAI22_X1 i_0_0_187 (.A1(n_0_0_353), .A2(n_0_0_319), .B1(shamt[0]), .B2(
      n_0_0_323), .ZN(Nb[14]));
   AOI22_X1 i_0_0_194 (.A1(shamt[1]), .A2(n_0_0_397), .B1(n_0_0_355), .B2(
      n_0_0_327), .ZN(n_0_0_319));
   OAI22_X1 i_0_0_195 (.A1(n_0_0_353), .A2(n_0_0_323), .B1(shamt[0]), .B2(
      n_0_0_326), .ZN(Nb[15]));
   AOI22_X1 i_0_0_196 (.A1(n_0_0_355), .A2(n_0_0_330), .B1(shamt[1]), .B2(
      n_0_0_324), .ZN(n_0_0_323));
   AOI22_X1 i_0_0_209 (.A1(n_0_0_70), .A2(n_0_0_337), .B1(shamt[2]), .B2(
      n_0_0_384), .ZN(n_0_0_324));
   OAI22_X1 i_0_0_210 (.A1(n_0_0_353), .A2(n_0_0_326), .B1(shamt[0]), .B2(
      n_0_0_329), .ZN(Nb[16]));
   AOI22_X1 i_0_0_211 (.A1(n_0_0_355), .A2(n_0_0_333), .B1(shamt[1]), .B2(
      n_0_0_327), .ZN(n_0_0_326));
   AOI22_X1 i_0_0_213 (.A1(n_0_0_70), .A2(n_0_0_340), .B1(shamt[2]), .B2(
      n_0_0_366), .ZN(n_0_0_327));
   OAI22_X1 i_0_0_214 (.A1(n_0_0_353), .A2(n_0_0_329), .B1(shamt[0]), .B2(
      n_0_0_332), .ZN(Nb[17]));
   AOI22_X1 i_0_0_216 (.A1(n_0_0_355), .A2(n_0_0_336), .B1(shamt[1]), .B2(
      n_0_0_330), .ZN(n_0_0_329));
   AOI22_X1 i_0_0_217 (.A1(n_0_0_70), .A2(n_0_0_343), .B1(shamt[2]), .B2(
      n_0_0_401), .ZN(n_0_0_330));
   OAI22_X1 i_0_0_218 (.A1(n_0_0_353), .A2(n_0_0_332), .B1(shamt[0]), .B2(
      n_0_0_335), .ZN(Nb[18]));
   AOI22_X1 i_0_0_219 (.A1(n_0_0_355), .A2(n_0_0_339), .B1(shamt[1]), .B2(
      n_0_0_333), .ZN(n_0_0_332));
   AOI22_X1 i_0_0_220 (.A1(n_0_0_70), .A2(n_0_0_346), .B1(shamt[2]), .B2(
      n_0_0_398), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_221 (.A1(n_0_0_353), .A2(n_0_0_335), .B1(shamt[0]), .B2(
      n_0_0_338), .ZN(Nb[19]));
   AOI22_X1 i_0_0_222 (.A1(shamt[1]), .A2(n_0_0_336), .B1(n_0_0_355), .B2(
      n_0_0_342), .ZN(n_0_0_335));
   OAI22_X1 i_0_0_223 (.A1(n_0_0_70), .A2(n_0_0_337), .B1(shamt[2]), .B2(
      n_0_0_374), .ZN(n_0_0_336));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_385), .A2(n_0_65), .B1(n_0_0_331), .B2(n_0_73), 
      .ZN(n_0_0_337));
   OAI22_X1 i_0_0_225 (.A1(n_0_0_353), .A2(n_0_0_338), .B1(shamt[0]), .B2(
      n_0_0_341), .ZN(Nb[20]));
   AOI22_X1 i_0_0_226 (.A1(n_0_0_355), .A2(n_0_0_345), .B1(shamt[1]), .B2(
      n_0_0_339), .ZN(n_0_0_338));
   OAI22_X1 i_0_0_227 (.A1(n_0_0_70), .A2(n_0_0_340), .B1(shamt[2]), .B2(
      n_0_0_363), .ZN(n_0_0_339));
   AOI22_X1 i_0_0_228 (.A1(n_0_0_385), .A2(n_0_66), .B1(n_0_0_331), .B2(n_0_74), 
      .ZN(n_0_0_340));
   OAI22_X1 i_0_0_229 (.A1(n_0_0_353), .A2(n_0_0_341), .B1(shamt[0]), .B2(
      n_0_0_344), .ZN(Nb[21]));
   AOI22_X1 i_0_0_230 (.A1(n_0_0_355), .A2(n_0_0_373), .B1(shamt[1]), .B2(
      n_0_0_342), .ZN(n_0_0_341));
   OAI22_X1 i_0_0_231 (.A1(n_0_0_70), .A2(n_0_0_343), .B1(shamt[2]), .B2(
      n_0_0_382), .ZN(n_0_0_342));
   AOI22_X1 i_0_0_232 (.A1(n_0_75), .A2(n_0_0_331), .B1(n_0_0_385), .B2(n_0_67), 
      .ZN(n_0_0_343));
   OAI22_X1 i_0_0_233 (.A1(n_0_0_353), .A2(n_0_0_344), .B1(shamt[0]), .B2(
      n_0_0_371), .ZN(Nb[22]));
   AOI22_X1 i_0_0_234 (.A1(shamt[1]), .A2(n_0_0_345), .B1(n_0_0_355), .B2(
      n_0_0_362), .ZN(n_0_0_344));
   OAI22_X1 i_0_0_235 (.A1(n_0_0_70), .A2(n_0_0_346), .B1(shamt[2]), .B2(
      n_0_0_352), .ZN(n_0_0_345));
   AOI22_X1 i_0_0_236 (.A1(n_0_0_331), .A2(n_0_76), .B1(n_0_0_385), .B2(n_0_68), 
      .ZN(n_0_0_346));
   OAI21_X1 i_0_0_237 (.A(n_0_0_347), .B1(n_0_0_353), .B2(n_0_0_371), .ZN(Nb[23]));
   OAI21_X1 i_0_0_238 (.A(n_0_0_348), .B1(n_0_0_355), .B2(n_0_0_362), .ZN(
      n_0_0_347));
   AOI21_X1 i_0_0_239 (.A(shamt[0]), .B1(n_0_0_355), .B2(n_0_0_349), .ZN(
      n_0_0_348));
   AOI22_X1 i_0_0_240 (.A1(n_0_0_360), .A2(n_0_0_350), .B1(shamt[2]), .B2(
      n_0_0_351), .ZN(n_0_0_349));
   AOI221_X1 i_0_0_241 (.A(shamt[2]), .B1(n_0_0_331), .B2(n_0_0_356), .C1(
      n_0_0_385), .C2(n_0_0_359), .ZN(n_0_0_350));
   INV_X1 i_0_0_242 (.A(n_0_0_352), .ZN(n_0_0_351));
   AOI222_X1 i_0_0_243 (.A1(n_0_0_331), .A2(n_0_80), .B1(n_0_0_388), .B2(n_0_64), 
      .C1(n_0_0_385), .C2(n_0_72), .ZN(n_0_0_352));
   INV_X1 i_0_0_244 (.A(n_0_0_354), .ZN(n_0_80));
   AOI22_X1 i_0_0_245 (.A1(n_0_10), .A2(n_0_0_37), .B1(n_0_41), .B2(n_0_0_36), 
      .ZN(n_0_0_354));
   INV_X1 i_0_0_246 (.A(n_0_0_356), .ZN(n_0_84));
   NAND2_X1 i_0_0_247 (.A1(n_0_0_37), .A2(n_0_0_46), .ZN(n_0_0_356));
   INV_X1 i_0_0_264 (.A(n_0_0_359), .ZN(n_0_76));
   AOI22_X1 i_0_0_265 (.A1(n_0_14), .A2(n_0_0_37), .B1(n_0_45), .B2(n_0_0_36), 
      .ZN(n_0_0_359));
   OAI21_X1 i_0_0_266 (.A(shamt[4]), .B1(shamt[3]), .B2(n_0_0_361), .ZN(
      n_0_0_360));
   AOI22_X1 i_0_0_267 (.A1(shamt[2]), .A2(n_0_0_363), .B1(n_0_0_70), .B2(
      n_0_0_367), .ZN(n_0_0_362));
   AOI222_X1 i_0_0_268 (.A1(n_0_0_331), .A2(n_0_78), .B1(n_0_0_385), .B2(n_0_70), 
      .C1(n_0_0_388), .C2(n_0_62), .ZN(n_0_0_363));
   INV_X1 i_0_0_269 (.A(n_0_0_365), .ZN(n_0_78));
   AOI22_X1 i_0_0_270 (.A1(n_0_12), .A2(n_0_0_37), .B1(n_0_43), .B2(n_0_0_36), 
      .ZN(n_0_0_365));
   AOI222_X1 i_0_0_271 (.A1(n_0_0_388), .A2(n_0_66), .B1(n_0_0_331), .B2(n_0_82), 
      .C1(n_0_0_385), .C2(n_0_74), .ZN(n_0_0_367));
   INV_X1 i_0_0_272 (.A(n_0_0_368), .ZN(n_0_82));
   AOI22_X1 i_0_0_273 (.A1(n_0_8), .A2(n_0_0_37), .B1(n_0_39), .B2(n_0_0_36), 
      .ZN(n_0_0_368));
   INV_X1 i_0_0_274 (.A(n_0_0_370), .ZN(n_0_74));
   OAI22_X1 i_0_0_275 (.A1(n_0_47), .A2(n_0_0_37), .B1(n_0_16), .B2(n_0_0_36), 
      .ZN(n_0_0_370));
   AOI21_X1 i_0_0_276 (.A(n_0_0_372), .B1(shamt[1]), .B2(n_0_0_373), .ZN(
      n_0_0_371));
   AOI221_X1 i_0_0_277 (.A(shamt[1]), .B1(n_0_0_70), .B2(n_0_0_386), .C1(
      shamt[2]), .C2(n_0_0_382), .ZN(n_0_0_372));
   AOI22_X1 i_0_0_278 (.A1(shamt[2]), .A2(n_0_0_374), .B1(n_0_0_70), .B2(
      n_0_0_378), .ZN(n_0_0_373));
   AOI222_X1 i_0_0_279 (.A1(n_0_0_331), .A2(n_0_77), .B1(n_0_0_385), .B2(n_0_69), 
      .C1(n_0_0_388), .C2(n_0_61), .ZN(n_0_0_374));
   INV_X1 i_0_0_280 (.A(n_0_0_376), .ZN(n_0_77));
   AOI22_X1 i_0_0_281 (.A1(n_0_13), .A2(n_0_0_37), .B1(n_0_44), .B2(n_0_0_36), 
      .ZN(n_0_0_376));
   AOI222_X1 i_0_0_282 (.A1(n_0_0_385), .A2(n_0_73), .B1(n_0_0_331), .B2(n_0_81), 
      .C1(n_0_0_388), .C2(n_0_65), .ZN(n_0_0_378));
   INV_X1 i_0_0_283 (.A(n_0_0_379), .ZN(n_0_81));
   AOI22_X1 i_0_0_284 (.A1(n_0_9), .A2(n_0_0_37), .B1(n_0_40), .B2(n_0_0_36), 
      .ZN(n_0_0_379));
   INV_X1 i_0_0_285 (.A(n_0_0_380), .ZN(n_0_73));
   OAI22_X1 i_0_0_286 (.A1(n_0_48), .A2(n_0_0_37), .B1(n_0_17), .B2(n_0_0_36), 
      .ZN(n_0_0_380));
   AOI222_X1 i_0_0_287 (.A1(n_0_0_388), .A2(n_0_63), .B1(n_0_0_331), .B2(n_0_79), 
      .C1(n_0_0_385), .C2(n_0_71), .ZN(n_0_0_382));
   INV_X1 i_0_0_288 (.A(n_0_0_383), .ZN(n_0_79));
   AOI22_X1 i_0_0_289 (.A1(n_0_11), .A2(n_0_0_37), .B1(n_0_42), .B2(n_0_0_36), 
      .ZN(n_0_0_383));
   AOI222_X1 i_0_0_290 (.A1(n_0_0_385), .A2(n_0_75), .B1(n_0_0_388), .B2(n_0_67), 
      .C1(n_0_0_331), .C2(n_0_83), .ZN(n_0_0_386));
   NOR2_X1 i_0_0_291 (.A1(n_0_0_394), .A2(shamt[3]), .ZN(n_0_0_388));
   INV_X1 i_0_0_292 (.A(n_0_0_389), .ZN(n_0_83));
   AOI22_X1 i_0_0_293 (.A1(n_0_7), .A2(n_0_0_37), .B1(n_0_38), .B2(n_0_0_36), 
      .ZN(n_0_0_389));
   INV_X1 i_0_0_294 (.A(n_0_0_391), .ZN(n_0_75));
   AOI22_X1 i_0_0_295 (.A1(n_0_15), .A2(n_0_0_37), .B1(n_0_46), .B2(n_0_0_36), 
      .ZN(n_0_0_391));
   INV_X1 i_0_0_296 (.A(mult_res[47]), .ZN(n_0_0_12));
   INV_X1 i_0_0_297 (.A(outA[0]), .ZN(n_0_0_35));
   NOR3_X1 i_0_0_298 (.A1(n_0_0_35), .A2(outA[1]), .A3(outA[2]), .ZN(n_0_0_36));
   INV_X1 i_0_0_299 (.A(n_0_0_36), .ZN(n_0_0_37));
   AOI22_X1 i_0_0_300 (.A1(n_0_0_37), .A2(n_0_35), .B1(n_0_0_36), .B2(n_0_5), 
      .ZN(n_0_0_38));
   XOR2_X1 i_0_0_348 (.A(n_0_0_38), .B(shamt[2]), .Z(n_0_0_39));
   INV_X1 i_0_0_349 (.A(b), .ZN(n_0_0_40));
   INV_X1 i_0_0_350 (.A(outB[0]), .ZN(n_0_0_41));
   NOR3_X1 i_0_0_351 (.A1(n_0_0_41), .A2(outB[1]), .A3(outB[2]), .ZN(n_0_0_45));
   INV_X1 i_0_0_352 (.A(n_0_0_45), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_353 (.A1(n_0_0_46), .A2(n_0_0_40), .ZN(n_0_0_47));
   AOI22_X1 i_0_0_354 (.A1(n_0_0_37), .A2(n_0_37), .B1(n_0_0_47), .B2(n_0_0_36), 
      .ZN(n_0_0_48));
   NAND2_X1 i_0_0_355 (.A1(n_0_0_48), .A2(shamt[0]), .ZN(n_0_0_49));
   OAI22_X1 i_0_0_356 (.A1(n_0_0_37), .A2(n_0_6), .B1(n_0_0_36), .B2(n_0_36), 
      .ZN(n_0_0_53));
   NAND2_X1 i_0_0_357 (.A1(n_0_0_53), .A2(shamt[1]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_358 (.A(n_0_0_54), .B1(n_0_0_53), .B2(shamt[1]), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_359 (.A(n_0_0_54), .B1(n_0_0_55), .B2(n_0_0_49), .ZN(n_0_0_56));
   AOI22_X1 i_0_0_360 (.A1(n_0_0_56), .A2(n_0_0_39), .B1(n_0_0_38), .B2(shamt[2]), 
      .ZN(n_0_0_60));
   OAI22_X1 i_0_0_361 (.A1(n_0_0_37), .A2(n_0_4), .B1(n_0_0_36), .B2(n_0_34), 
      .ZN(n_0_0_61));
   OR2_X1 i_0_0_362 (.A1(n_0_0_61), .A2(shamt[3]), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_363 (.A1(n_0_0_61), .A2(shamt[3]), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_364 (.A1(n_0_0_62), .A2(n_0_0_63), .ZN(n_0_0_68));
   XNOR2_X1 i_0_0_365 (.A(n_0_0_60), .B(n_0_0_68), .ZN(n_0_0_69));
   INV_X1 i_0_0_366 (.A(shamt[2]), .ZN(n_0_0_70));
   AOI22_X1 i_0_0_367 (.A1(mult_res[23]), .A2(n_0_0_93), .B1(n_0_0_235), 
      .B2(n_0_0_76), .ZN(n_0_0_75));
   AOI21_X1 i_0_0_368 (.A(n_0_0_77), .B1(E_sum[0]), .B2(n_0_0_94), .ZN(n_0_0_76));
   AOI221_X1 i_0_0_369 (.A(E_sum[0]), .B1(n_0_0_234), .B2(n_0_0_201), .C1(
      n_0_0_231), .C2(n_0_0_84), .ZN(n_0_0_77));
   AOI22_X1 i_0_0_370 (.A1(n_0_0_219), .A2(n_0_0_85), .B1(n_0_0_218), .B2(
      n_0_0_210), .ZN(n_0_0_84));
   AOI22_X1 i_0_0_371 (.A1(n_0_0_216), .A2(n_0_0_86), .B1(mult_res[31]), 
      .B2(n_0_0_213), .ZN(n_0_0_85));
   INV_X1 i_0_0_372 (.A(n_0_0_92), .ZN(n_0_0_86));
   AOI22_X1 i_0_0_373 (.A1(mult_res[23]), .A2(n_0_0_215), .B1(mult_res[39]), 
      .B2(n_0_0_214), .ZN(n_0_0_92));
   NOR3_X1 i_0_0_374 (.A1(n_0_0_248), .A2(n_0_0_242), .A3(mult_res[47]), 
      .ZN(n_0_0_93));
   OAI22_X1 i_0_0_375 (.A1(n_0_0_234), .A2(n_0_0_148), .B1(n_0_0_231), .B2(
      n_0_0_191), .ZN(n_0_0_94));
   AOI22_X1 i_0_0_376 (.A1(n_0_0_219), .A2(n_0_0_183), .B1(n_0_0_218), .B2(
      n_0_0_198), .ZN(n_0_0_148));
   AOI22_X1 i_0_0_377 (.A1(n_0_0_216), .A2(n_0_0_187), .B1(mult_res[32]), 
      .B2(n_0_0_213), .ZN(n_0_0_183));
   INV_X1 i_0_0_378 (.A(n_0_0_188), .ZN(n_0_0_187));
   OAI22_X1 i_0_0_379 (.A1(mult_res[24]), .A2(n_0_0_214), .B1(mult_res[40]), 
      .B2(n_0_0_215), .ZN(n_0_0_188));
   OAI22_X1 i_0_0_380 (.A1(n_0_0_218), .A2(n_0_0_192), .B1(n_0_0_219), .B2(
      n_0_0_195), .ZN(n_0_0_191));
   AOI22_X1 i_0_0_381 (.A1(mult_res[34]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_193), .ZN(n_0_0_192));
   INV_X1 i_0_0_382 (.A(n_0_0_194), .ZN(n_0_0_193));
   AOI22_X1 i_0_0_383 (.A1(mult_res[42]), .A2(n_0_0_214), .B1(mult_res[26]), 
      .B2(n_0_0_215), .ZN(n_0_0_194));
   AOI22_X1 i_0_0_384 (.A1(mult_res[38]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_196), .ZN(n_0_0_195));
   INV_X1 i_0_0_385 (.A(n_0_0_197), .ZN(n_0_0_196));
   OAI22_X1 i_0_0_386 (.A1(mult_res[46]), .A2(n_0_0_215), .B1(mult_res[30]), 
      .B2(n_0_0_214), .ZN(n_0_0_197));
   AOI22_X1 i_0_0_387 (.A1(mult_res[36]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_199), .ZN(n_0_0_198));
   INV_X1 i_0_0_388 (.A(n_0_0_200), .ZN(n_0_0_199));
   OAI22_X1 i_0_0_389 (.A1(mult_res[44]), .A2(n_0_0_215), .B1(mult_res[28]), 
      .B2(n_0_0_214), .ZN(n_0_0_200));
   OAI22_X1 i_0_0_390 (.A1(n_0_0_218), .A2(n_0_0_202), .B1(n_0_0_219), .B2(
      n_0_0_206), .ZN(n_0_0_201));
   AOI22_X1 i_0_0_391 (.A1(mult_res[33]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_203), .ZN(n_0_0_202));
   INV_X1 i_0_0_392 (.A(n_0_0_204), .ZN(n_0_0_203));
   AOI22_X1 i_0_0_393 (.A1(mult_res[41]), .A2(n_0_0_214), .B1(mult_res[25]), 
      .B2(n_0_0_215), .ZN(n_0_0_204));
   AOI22_X1 i_0_0_394 (.A1(mult_res[37]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_207), .ZN(n_0_0_206));
   INV_X1 i_0_0_395 (.A(n_0_0_209), .ZN(n_0_0_207));
   OAI22_X1 i_0_0_396 (.A1(mult_res[29]), .A2(n_0_0_214), .B1(mult_res[45]), 
      .B2(n_0_0_215), .ZN(n_0_0_209));
   AOI22_X1 i_0_0_397 (.A1(mult_res[35]), .A2(n_0_0_213), .B1(n_0_0_216), 
      .B2(n_0_0_211), .ZN(n_0_0_210));
   INV_X1 i_0_0_398 (.A(n_0_0_212), .ZN(n_0_0_211));
   OAI22_X1 i_0_0_399 (.A1(mult_res[27]), .A2(n_0_0_214), .B1(mult_res[43]), 
      .B2(n_0_0_215), .ZN(n_0_0_212));
   NOR2_X1 i_0_0_400 (.A1(n_0_0_216), .A2(n_0_0_214), .ZN(n_0_0_213));
   INV_X1 i_0_0_401 (.A(n_0_0_215), .ZN(n_0_0_214));
   OAI21_X1 i_0_0_402 (.A(n_0_0_238), .B1(n_0_0_305), .B2(n_0_0_239), .ZN(
      n_0_0_215));
   INV_X1 i_0_0_403 (.A(n_0_0_217), .ZN(n_0_0_216));
   AOI21_X1 i_0_0_404 (.A(n_0_0_239), .B1(E_sum[3]), .B2(n_0_0_240), .ZN(
      n_0_0_217));
   INV_X1 i_0_0_405 (.A(n_0_0_219), .ZN(n_0_0_218));
   OAI21_X1 i_0_0_406 (.A(n_0_0_240), .B1(n_0_0_304), .B2(n_0_0_241), .ZN(
      n_0_0_219));
   INV_X1 i_0_0_407 (.A(n_0_0_234), .ZN(n_0_0_231));
   OAI22_X1 i_0_0_408 (.A1(n_0_0_303), .A2(E_sum[0]), .B1(E_sum[1]), .B2(
      n_0_0_302), .ZN(n_0_0_234));
   AOI211_X1 i_0_0_409 (.A(n_0_0_243), .B(n_0_0_248), .C1(n_0_0_237), .C2(
      n_0_0_236), .ZN(n_0_0_235));
   OR4_X1 i_0_0_410 (.A1(E_sum[6]), .A2(n_0_0_238), .A3(E_sum[5]), .A4(n_0_0_306), 
      .ZN(n_0_0_236));
   NAND4_X1 i_0_0_411 (.A1(E_sum[6]), .A2(n_0_0_238), .A3(E_sum[5]), .A4(
      n_0_0_306), .ZN(n_0_0_237));
   NAND2_X1 i_0_0_412 (.A1(n_0_0_305), .A2(n_0_0_239), .ZN(n_0_0_238));
   NOR2_X1 i_0_0_413 (.A1(E_sum[3]), .A2(n_0_0_240), .ZN(n_0_0_239));
   NAND2_X1 i_0_0_414 (.A1(n_0_0_304), .A2(n_0_0_241), .ZN(n_0_0_240));
   NOR2_X1 i_0_0_415 (.A1(E_sum[1]), .A2(E_sum[0]), .ZN(n_0_0_241));
   INV_X1 i_0_0_416 (.A(n_0_0_243), .ZN(n_0_0_242));
   AOI21_X1 i_0_0_417 (.A(n_0_0_247), .B1(n_0_0_246), .B2(n_0_0_244), .ZN(
      n_0_0_243));
   AND2_X1 i_0_0_418 (.A1(n_0_0_255), .A2(n_0_0_245), .ZN(n_0_0_244));
   NOR4_X1 i_0_0_419 (.A1(n_0_0_302), .A2(n_0_0_13), .A3(n_0_0_14), .A4(n_0_0_15), 
      .ZN(n_0_0_245));
   NOR4_X1 i_0_0_420 (.A1(n_0_0_17), .A2(n_0_0_16), .A3(n_0_0_18), .A4(n_0_0_253), 
      .ZN(n_0_0_246));
   OAI21_X1 i_0_0_421 (.A(n_0_0_257), .B1(E_sum[8]), .B2(n_0_0_255), .ZN(
      n_0_0_247));
   NAND3_X1 i_0_0_422 (.A1(n_0_0_257), .A2(n_0_0_249), .A3(enable), .ZN(
      n_0_0_248));
   AOI21_X1 i_0_0_423 (.A(n_0_0_250), .B1(E_sum[8]), .B2(n_0_0_255), .ZN(
      n_0_0_249));
   NOR3_X1 i_0_0_424 (.A1(n_0_0_252), .A2(n_0_0_251), .A3(n_0_0_254), .ZN(
      n_0_0_250));
   NAND4_X1 i_0_0_425 (.A1(n_0_0_17), .A2(n_0_0_16), .A3(n_0_0_302), .A4(
      n_0_0_18), .ZN(n_0_0_251));
   NAND3_X1 i_0_0_426 (.A1(n_0_0_15), .A2(n_0_0_14), .A3(n_0_0_13), .ZN(
      n_0_0_252));
   INV_X1 i_0_0_427 (.A(n_0_0_254), .ZN(n_0_0_253));
   AOI21_X1 i_0_0_428 (.A(E_sum[8]), .B1(E_sum[7]), .B2(n_0_0_28), .ZN(n_0_0_254));
   INV_X1 i_0_0_429 (.A(n_0_0_256), .ZN(n_0_0_255));
   NOR2_X1 i_0_0_430 (.A1(E_sum[7]), .A2(n_0_0_28), .ZN(n_0_0_256));
   NAND2_X1 i_0_0_431 (.A1(n_0_0_259), .A2(n_0_0_258), .ZN(n_0_0_257));
   AOI22_X1 i_0_0_432 (.A1(n_0_0), .A2(n_0_0_36), .B1(n_0_0_37), .B2(n_0_30), 
      .ZN(n_0_0_258));
   INV_X1 i_0_0_433 (.A(n_0_0_260), .ZN(n_0_0_259));
   NAND2_X1 i_0_0_434 (.A1(n_0_0_262), .A2(n_0_0_261), .ZN(n_0_0_260));
   AOI22_X1 i_0_0_435 (.A1(n_0_1), .A2(n_0_0_36), .B1(n_0_0_37), .B2(n_0_31), 
      .ZN(n_0_0_261));
   INV_X1 i_0_0_436 (.A(n_0_0_263), .ZN(n_0_0_262));
   NAND2_X1 i_0_0_437 (.A1(n_0_0_294), .A2(n_0_0_265), .ZN(n_0_0_263));
   AOI22_X1 i_0_0_438 (.A1(n_0_2), .A2(n_0_0_36), .B1(n_0_0_37), .B2(n_0_32), 
      .ZN(n_0_0_265));
   AOI21_X1 i_0_0_439 (.A(n_0_0_299), .B1(n_0_0_296), .B2(n_0_0_295), .ZN(
      n_0_0_294));
   NAND2_X1 i_0_0_440 (.A1(shamt[4]), .A2(n_0_0_301), .ZN(n_0_0_295));
   NAND2_X1 i_0_0_441 (.A1(n_0_0_62), .A2(n_0_0_298), .ZN(n_0_0_296));
   NAND2_X1 i_0_0_442 (.A1(n_0_0_60), .A2(n_0_0_63), .ZN(n_0_0_298));
   NOR2_X1 i_0_0_443 (.A1(shamt[4]), .A2(n_0_0_301), .ZN(n_0_0_299));
   OAI22_X1 i_0_0_444 (.A1(n_0_33), .A2(n_0_0_36), .B1(n_0_3), .B2(n_0_0_37), 
      .ZN(n_0_0_301));
   INV_X1 i_0_0_445 (.A(E_sum[0]), .ZN(n_0_0_302));
   INV_X1 i_0_0_446 (.A(E_sum[1]), .ZN(n_0_0_303));
   INV_X1 i_0_0_447 (.A(E_sum[2]), .ZN(n_0_0_304));
   INV_X1 i_0_0_448 (.A(E_sum[4]), .ZN(n_0_0_305));
   INV_X1 i_0_0_449 (.A(E_sum[7]), .ZN(n_0_0_306));
   OAI22_X1 i_0_0_450 (.A1(n_0_0_309), .A2(n_0_0_307), .B1(enable), .B2(
      n_0_0_308), .ZN(res[31]));
   XNOR2_X1 i_0_0_451 (.A(Sa), .B(Sb), .ZN(n_0_0_307));
   INV_X1 i_0_0_452 (.A(special_res[31]), .ZN(n_0_0_308));
   INV_X1 i_0_0_453 (.A(enable), .ZN(n_0_0_309));
   AOI22_X1 i_0_0_454 (.A1(n_0_0_353), .A2(n_0_0_310), .B1(shamt[0]), .B2(
      n_0_0_315), .ZN(Nb[5]));
   AOI22_X1 i_0_0_455 (.A1(n_0_0_355), .A2(n_0_0_312), .B1(n_0_0_317), .B2(
      n_0_64), .ZN(n_0_0_310));
   INV_X1 i_0_0_456 (.A(n_0_0_311), .ZN(n_0_64));
   OAI22_X1 i_0_0_457 (.A1(n_0_57), .A2(n_0_0_37), .B1(n_0_26), .B2(n_0_0_36), 
      .ZN(n_0_0_311));
   OAI22_X1 i_0_0_458 (.A1(n_0_0_325), .A2(n_0_0_314), .B1(n_0_0_321), .B2(
      n_0_0_313), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_459 (.A1(n_0_55), .A2(n_0_0_37), .B1(n_0_24), .B2(n_0_0_36), 
      .ZN(n_0_0_313));
   INV_X1 i_0_0_460 (.A(n_0_0_314), .ZN(n_0_62));
   OAI22_X1 i_0_0_461 (.A1(n_0_59), .A2(n_0_0_37), .B1(n_0_28), .B2(n_0_0_36), 
      .ZN(n_0_0_314));
   AOI22_X1 i_0_0_462 (.A1(n_0_0_355), .A2(n_0_0_320), .B1(n_0_63), .B2(
      n_0_0_317), .ZN(n_0_0_315));
   NOR2_X1 i_0_0_463 (.A1(n_0_0_355), .A2(n_0_0_321), .ZN(n_0_0_317));
   INV_X1 i_0_0_464 (.A(n_0_0_318), .ZN(n_0_63));
   OAI22_X1 i_0_0_465 (.A1(n_0_58), .A2(n_0_0_37), .B1(n_0_27), .B2(n_0_0_36), 
      .ZN(n_0_0_318));
   OAI22_X1 i_0_0_466 (.A1(n_0_0_334), .A2(n_0_0_325), .B1(n_0_0_322), .B2(
      n_0_0_321), .ZN(n_0_0_320));
   NAND2_X1 i_0_0_467 (.A1(n_0_0_70), .A2(n_0_0_331), .ZN(n_0_0_321));
   OAI22_X1 i_0_0_468 (.A1(n_0_56), .A2(n_0_0_37), .B1(n_0_25), .B2(n_0_0_36), 
      .ZN(n_0_0_322));
   INV_X1 i_0_0_469 (.A(n_0_0_328), .ZN(n_0_0_325));
   NOR3_X1 i_0_0_470 (.A1(shamt[4]), .A2(shamt[3]), .A3(n_0_0_70), .ZN(n_0_0_328));
   NOR2_X1 i_0_0_471 (.A1(shamt[4]), .A2(shamt[3]), .ZN(n_0_0_331));
   INV_X1 i_0_0_472 (.A(n_0_0_334), .ZN(n_0_61));
   OAI22_X1 i_0_0_473 (.A1(n_0_60), .A2(n_0_0_37), .B1(n_0_29), .B2(n_0_0_36), 
      .ZN(n_0_0_334));
   INV_X1 i_0_0_474 (.A(shamt[0]), .ZN(n_0_0_353));
   INV_X1 i_0_0_475 (.A(shamt[1]), .ZN(n_0_0_355));
   OAI22_X1 i_0_0_476 (.A1(shamt[0]), .A2(n_0_0_357), .B1(n_0_0_353), .B2(
      n_0_0_369), .ZN(Nb[9]));
   AOI22_X1 i_0_0_477 (.A1(n_0_0_355), .A2(n_0_0_364), .B1(shamt[1]), .B2(
      n_0_0_358), .ZN(n_0_0_357));
   OAI22_X1 i_0_0_478 (.A1(n_0_0_395), .A2(n_0_0_393), .B1(n_0_0_321), .B2(
      n_0_0_361), .ZN(n_0_0_358));
   OAI22_X1 i_0_0_479 (.A1(n_0_22), .A2(n_0_0_36), .B1(n_0_0_37), .B2(n_0_53), 
      .ZN(n_0_0_361));
   OAI22_X1 i_0_0_480 (.A1(n_0_0_395), .A2(n_0_0_313), .B1(shamt[2]), .B2(
      n_0_0_366), .ZN(n_0_0_364));
   AOI22_X1 i_0_0_481 (.A1(n_0_0_331), .A2(n_0_70), .B1(n_0_62), .B2(n_0_0_385), 
      .ZN(n_0_0_366));
   AOI22_X1 i_0_0_482 (.A1(n_0_0_355), .A2(n_0_0_381), .B1(shamt[1]), .B2(
      n_0_0_375), .ZN(n_0_0_369));
   OAI22_X1 i_0_0_483 (.A1(n_0_0_395), .A2(n_0_0_392), .B1(n_0_0_321), .B2(
      n_0_0_377), .ZN(n_0_0_375));
   OAI22_X1 i_0_0_484 (.A1(n_0_23), .A2(n_0_0_36), .B1(n_0_0_37), .B2(n_0_54), 
      .ZN(n_0_0_377));
   OAI22_X1 i_0_0_485 (.A1(n_0_0_322), .A2(n_0_0_395), .B1(shamt[2]), .B2(
      n_0_0_384), .ZN(n_0_0_381));
   AOI22_X1 i_0_0_486 (.A1(n_0_0_331), .A2(n_0_69), .B1(n_0_61), .B2(n_0_0_385), 
      .ZN(n_0_0_384));
   AND2_X1 i_0_0_487 (.A1(n_0_0_394), .A2(shamt[3]), .ZN(n_0_0_385));
   INV_X1 i_0_0_488 (.A(n_0_0_387), .ZN(n_0_69));
   AOI22_X1 i_0_0_489 (.A1(n_0_21), .A2(n_0_0_37), .B1(n_0_52), .B2(n_0_0_36), 
      .ZN(n_0_0_387));
   INV_X1 i_0_0_490 (.A(n_0_0_390), .ZN(n_0_70));
   AOI22_X1 i_0_0_491 (.A1(n_0_20), .A2(n_0_0_37), .B1(n_0_51), .B2(n_0_0_36), 
      .ZN(n_0_0_390));
   INV_X1 i_0_0_492 (.A(n_0_0_313), .ZN(n_0_66));
   INV_X1 i_0_0_493 (.A(n_0_63), .ZN(n_0_0_392));
   INV_X1 i_0_0_494 (.A(n_0_64), .ZN(n_0_0_393));
   INV_X1 i_0_0_495 (.A(shamt[4]), .ZN(n_0_0_394));
   INV_X1 i_0_0_496 (.A(n_0_0_328), .ZN(n_0_0_395));
   INV_X1 i_0_0_497 (.A(n_0_0_322), .ZN(n_0_65));
   OAI22_X1 i_0_0_498 (.A1(shamt[0]), .A2(n_0_0_396), .B1(n_0_0_353), .B2(
      n_0_0_399), .ZN(Nb[11]));
   AOI22_X1 i_0_0_499 (.A1(shamt[1]), .A2(n_0_0_364), .B1(n_0_0_355), .B2(
      n_0_0_397), .ZN(n_0_0_396));
   OAI22_X1 i_0_0_500 (.A1(n_0_0_404), .A2(n_0_0_361), .B1(shamt[2]), .B2(
      n_0_0_398), .ZN(n_0_0_397));
   AOI22_X1 i_0_0_501 (.A1(n_0_0_331), .A2(n_0_72), .B1(n_0_0_385), .B2(n_0_64), 
      .ZN(n_0_0_398));
   AOI22_X1 i_0_0_502 (.A1(shamt[1]), .A2(n_0_0_381), .B1(n_0_0_355), .B2(
      n_0_0_400), .ZN(n_0_0_399));
   OAI22_X1 i_0_0_503 (.A1(n_0_0_377), .A2(n_0_0_404), .B1(shamt[2]), .B2(
      n_0_0_401), .ZN(n_0_0_400));
   AOI22_X1 i_0_0_504 (.A1(n_0_0_331), .A2(n_0_71), .B1(n_0_0_385), .B2(n_0_63), 
      .ZN(n_0_0_401));
   INV_X1 i_0_0_505 (.A(n_0_0_402), .ZN(n_0_71));
   AOI22_X1 i_0_0_506 (.A1(n_0_19), .A2(n_0_0_37), .B1(n_0_50), .B2(n_0_0_36), 
      .ZN(n_0_0_402));
   INV_X1 i_0_0_507 (.A(n_0_0_403), .ZN(n_0_72));
   AOI22_X1 i_0_0_508 (.A1(n_0_18), .A2(n_0_0_37), .B1(n_0_49), .B2(n_0_0_36), 
      .ZN(n_0_0_403));
   INV_X1 i_0_0_509 (.A(n_0_0_361), .ZN(n_0_68));
   INV_X1 i_0_0_510 (.A(n_0_0_328), .ZN(n_0_0_404));
   INV_X1 i_0_0_511 (.A(n_0_0_377), .ZN(n_0_67));
endmodule
