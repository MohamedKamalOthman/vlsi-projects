/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed Nov  2 22:05:53 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 348179448 */

module halfAdder__0_11(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_12(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   halfAdder__0_11 h1 (.in1(x), .in2(y), .cout(cout), .sum(sum));
endmodule

module halfAdder__0_19(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_16(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_20(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_19 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_16 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_27(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_24(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_28(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_27 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_24 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_35(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_32(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_36(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_35 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_32 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_43(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_40(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_44(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_43 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_40 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_51(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_48(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_52(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_51 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_48 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_59(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_56(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_60(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_59 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_56 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_67(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_64(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_68(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_67 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_64 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_75(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_72(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_76(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_75 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_72 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_83(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_80(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_84(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_83 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_80 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_91(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_88(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_92(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_91 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_88 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_99(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_96(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_100(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_99 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_96 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_107(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_104(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_108(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_107 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_104 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_115(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_112(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_116(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_115 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_112 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_123(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_120(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_124(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_123 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_120 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_131(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_128(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_132(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_131 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_128 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_139(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_136(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_140(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_139 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_136 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_147(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_144(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_148(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_147 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_144 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_155(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_152(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_156(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_155 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_152 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_163(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_160(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_164(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_163 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_160 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_171(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_168(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_172(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_171 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_168 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_179(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_176(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_180(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_179 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_176 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_187(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_184(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_188(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_187 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_184 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_195(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_192(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_196(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_195 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_192 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_203(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_200(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_204(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_203 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_200 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_211(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_208(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_212(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_211 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_208 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_219(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_216(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_220(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_219 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_216 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_227(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_224(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_228(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_227 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_224 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_235(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_232(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_236(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_235 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_232 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_243(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_240(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_244(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_243 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_240 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_251(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder__0_248(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder__0_252(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_251 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder__0_248 h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), 
      .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module halfAdder__0_4(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module halfAdder(in1, in2, cout, sum);
   input in1;
   input in2;
   output cout;
   output sum;

   AND2_X1 i_0_0 (.A1(in1), .A2(in2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1), .B(in2), .Z(sum));
endmodule

module fullAdder(cin, x, y, cout, sum);
   input cin;
   input x;
   input y;
   output cout;
   output sum;

   wire dummySum1;
   wire dummyCarry1;
   wire dummyCarry2;

   halfAdder__0_4 h1 (.in1(x), .in2(y), .cout(dummyCarry1), .sum(dummySum1));
   halfAdder h2d (.in1(dummySum1), .in2(cin), .cout(dummyCarry2), .sum(sum));
   OR2_X1 i_0_0 (.A1(dummyCarry1), .A2(dummyCarry2), .ZN(cout));
endmodule

module CarryRippleAdder(add1_i, add2_i, sum_o, carry_o);
   input [31:0]add1_i;
   input [31:0]add2_i;
   output [31:0]sum_o;
   output carry_o;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;

   fullAdder__0_12 genblk1_0_fa_inst (.cin(), .x(add1_i[0]), .y(add2_i[0]), 
      .cout(n_0_0), .sum(sum_o[0]));
   fullAdder__0_20 genblk1_1_fa_inst (.cin(n_0_0), .x(add1_i[1]), .y(add2_i[1]), 
      .cout(n_0_1), .sum(sum_o[1]));
   fullAdder__0_28 genblk1_2_fa_inst (.cin(n_0_1), .x(add1_i[2]), .y(add2_i[2]), 
      .cout(n_0_2), .sum(sum_o[2]));
   fullAdder__0_36 genblk1_3_fa_inst (.cin(n_0_2), .x(add1_i[3]), .y(add2_i[3]), 
      .cout(n_0_3), .sum(sum_o[3]));
   fullAdder__0_44 genblk1_4_fa_inst (.cin(n_0_3), .x(add1_i[4]), .y(add2_i[4]), 
      .cout(n_0_4), .sum(sum_o[4]));
   fullAdder__0_52 genblk1_5_fa_inst (.cin(n_0_4), .x(add1_i[5]), .y(add2_i[5]), 
      .cout(n_0_5), .sum(sum_o[5]));
   fullAdder__0_60 genblk1_6_fa_inst (.cin(n_0_5), .x(add1_i[6]), .y(add2_i[6]), 
      .cout(n_0_6), .sum(sum_o[6]));
   fullAdder__0_68 genblk1_7_fa_inst (.cin(n_0_6), .x(add1_i[7]), .y(add2_i[7]), 
      .cout(n_0_7), .sum(sum_o[7]));
   fullAdder__0_76 genblk1_8_fa_inst (.cin(n_0_7), .x(add1_i[8]), .y(add2_i[8]), 
      .cout(n_0_8), .sum(sum_o[8]));
   fullAdder__0_84 genblk1_9_fa_inst (.cin(n_0_8), .x(add1_i[9]), .y(add2_i[9]), 
      .cout(n_0_9), .sum(sum_o[9]));
   fullAdder__0_92 genblk1_10_fa_inst (.cin(n_0_9), .x(add1_i[10]), .y(
      add2_i[10]), .cout(n_0_10), .sum(sum_o[10]));
   fullAdder__0_100 genblk1_11_fa_inst (.cin(n_0_10), .x(add1_i[11]), .y(
      add2_i[11]), .cout(n_0_11), .sum(sum_o[11]));
   fullAdder__0_108 genblk1_12_fa_inst (.cin(n_0_11), .x(add1_i[12]), .y(
      add2_i[12]), .cout(n_0_12), .sum(sum_o[12]));
   fullAdder__0_116 genblk1_13_fa_inst (.cin(n_0_12), .x(add1_i[13]), .y(
      add2_i[13]), .cout(n_0_13), .sum(sum_o[13]));
   fullAdder__0_124 genblk1_14_fa_inst (.cin(n_0_13), .x(add1_i[14]), .y(
      add2_i[14]), .cout(n_0_14), .sum(sum_o[14]));
   fullAdder__0_132 genblk1_15_fa_inst (.cin(n_0_14), .x(add1_i[15]), .y(
      add2_i[15]), .cout(n_0_15), .sum(sum_o[15]));
   fullAdder__0_140 genblk1_16_fa_inst (.cin(n_0_15), .x(add1_i[16]), .y(
      add2_i[16]), .cout(n_0_16), .sum(sum_o[16]));
   fullAdder__0_148 genblk1_17_fa_inst (.cin(n_0_16), .x(add1_i[17]), .y(
      add2_i[17]), .cout(n_0_17), .sum(sum_o[17]));
   fullAdder__0_156 genblk1_18_fa_inst (.cin(n_0_17), .x(add1_i[18]), .y(
      add2_i[18]), .cout(n_0_18), .sum(sum_o[18]));
   fullAdder__0_164 genblk1_19_fa_inst (.cin(n_0_18), .x(add1_i[19]), .y(
      add2_i[19]), .cout(n_0_19), .sum(sum_o[19]));
   fullAdder__0_172 genblk1_20_fa_inst (.cin(n_0_19), .x(add1_i[20]), .y(
      add2_i[20]), .cout(n_0_20), .sum(sum_o[20]));
   fullAdder__0_180 genblk1_21_fa_inst (.cin(n_0_20), .x(add1_i[21]), .y(
      add2_i[21]), .cout(n_0_21), .sum(sum_o[21]));
   fullAdder__0_188 genblk1_22_fa_inst (.cin(n_0_21), .x(add1_i[22]), .y(
      add2_i[22]), .cout(n_0_22), .sum(sum_o[22]));
   fullAdder__0_196 genblk1_23_fa_inst (.cin(n_0_22), .x(add1_i[23]), .y(
      add2_i[23]), .cout(n_0_23), .sum(sum_o[23]));
   fullAdder__0_204 genblk1_24_fa_inst (.cin(n_0_23), .x(add1_i[24]), .y(
      add2_i[24]), .cout(n_0_24), .sum(sum_o[24]));
   fullAdder__0_212 genblk1_25_fa_inst (.cin(n_0_24), .x(add1_i[25]), .y(
      add2_i[25]), .cout(n_0_25), .sum(sum_o[25]));
   fullAdder__0_220 genblk1_26_fa_inst (.cin(n_0_25), .x(add1_i[26]), .y(
      add2_i[26]), .cout(n_0_26), .sum(sum_o[26]));
   fullAdder__0_228 genblk1_27_fa_inst (.cin(n_0_26), .x(add1_i[27]), .y(
      add2_i[27]), .cout(n_0_27), .sum(sum_o[27]));
   fullAdder__0_236 genblk1_28_fa_inst (.cin(n_0_27), .x(add1_i[28]), .y(
      add2_i[28]), .cout(n_0_28), .sum(sum_o[28]));
   fullAdder__0_244 genblk1_29_fa_inst (.cin(n_0_28), .x(add1_i[29]), .y(
      add2_i[29]), .cout(n_0_29), .sum(sum_o[29]));
   fullAdder__0_252 genblk1_30_fa_inst (.cin(n_0_29), .x(add1_i[30]), .y(
      add2_i[30]), .cout(n_0_30), .sum(sum_o[30]));
   fullAdder genblk1_31_fa_inst (.cin(n_0_30), .x(add1_i[31]), .y(add2_i[31]), 
      .cout(carry_o), .sum(sum_o[31]));
endmodule
