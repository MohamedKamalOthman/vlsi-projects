/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Mon Dec 26 10:55:55 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2218885896 */

module datapath(A, p_0, M_temp);
   input [31:0]A;
   output [31:0]p_0;
   input [31:0]M_temp;

   INV_X1 i_0 (.A(A[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(M_temp[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(M_temp[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(A[1]), .B(M_temp[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(A[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(M_temp[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(M_temp[2]), .B(A[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(M_temp[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(A[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(A[3]), .B(M_temp[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(A[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(M_temp[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(M_temp[4]), .B(A[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(M_temp[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(A[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(A[5]), .B(M_temp[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(A[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(M_temp[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(M_temp[6]), .B(A[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(M_temp[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(A[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(A[7]), .B(M_temp[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(A[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(M_temp[7]), .ZN(n_23));
   XOR2_X1 i_32 (.A(M_temp[8]), .B(A[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_0[8]));
   INV_X1 i_34 (.A(M_temp[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(A[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(A[9]), .B(M_temp[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_0[9]));
   INV_X1 i_38 (.A(A[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(M_temp[9]), .ZN(n_29));
   XOR2_X1 i_40 (.A(M_temp[10]), .B(A[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_0[10]));
   INV_X1 i_42 (.A(M_temp[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(A[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(A[11]), .B(M_temp[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_0[11]));
   INV_X1 i_46 (.A(A[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(M_temp[11]), .ZN(n_35));
   XOR2_X1 i_48 (.A(M_temp[12]), .B(A[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_0[12]));
   INV_X1 i_50 (.A(M_temp[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(A[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(A[13]), .B(M_temp[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_0[13]));
   INV_X1 i_54 (.A(A[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(M_temp[13]), .ZN(n_41));
   XOR2_X1 i_56 (.A(M_temp[14]), .B(A[14]), .Z(n_42));
   XNOR2_X1 i_57 (.A(n_41), .B(n_42), .ZN(p_0[14]));
   INV_X1 i_58 (.A(M_temp[14]), .ZN(n_43));
   OAI22_X1 i_59 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(A[14]), .ZN(n_44));
   XNOR2_X1 i_60 (.A(A[15]), .B(M_temp[15]), .ZN(n_45));
   XNOR2_X1 i_61 (.A(n_44), .B(n_45), .ZN(p_0[15]));
   INV_X1 i_62 (.A(A[15]), .ZN(n_46));
   AOI22_X1 i_63 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(M_temp[15]), .ZN(n_47));
   XOR2_X1 i_64 (.A(M_temp[16]), .B(A[16]), .Z(n_48));
   XNOR2_X1 i_65 (.A(n_47), .B(n_48), .ZN(p_0[16]));
   INV_X1 i_66 (.A(M_temp[16]), .ZN(n_49));
   OAI22_X1 i_67 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(A[16]), .ZN(n_50));
   XNOR2_X1 i_68 (.A(A[17]), .B(M_temp[17]), .ZN(n_51));
   XNOR2_X1 i_69 (.A(n_50), .B(n_51), .ZN(p_0[17]));
   INV_X1 i_70 (.A(A[17]), .ZN(n_52));
   AOI22_X1 i_71 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(M_temp[17]), .ZN(n_53));
   XOR2_X1 i_72 (.A(M_temp[18]), .B(A[18]), .Z(n_54));
   XNOR2_X1 i_73 (.A(n_53), .B(n_54), .ZN(p_0[18]));
   INV_X1 i_74 (.A(M_temp[18]), .ZN(n_55));
   OAI22_X1 i_75 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(A[18]), .ZN(n_56));
   XNOR2_X1 i_76 (.A(A[19]), .B(M_temp[19]), .ZN(n_57));
   XNOR2_X1 i_77 (.A(n_56), .B(n_57), .ZN(p_0[19]));
   INV_X1 i_78 (.A(A[19]), .ZN(n_58));
   AOI22_X1 i_79 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(M_temp[19]), .ZN(n_59));
   XOR2_X1 i_80 (.A(M_temp[20]), .B(A[20]), .Z(n_60));
   XNOR2_X1 i_81 (.A(n_59), .B(n_60), .ZN(p_0[20]));
   INV_X1 i_82 (.A(M_temp[20]), .ZN(n_61));
   OAI22_X1 i_83 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(A[20]), .ZN(n_62));
   XNOR2_X1 i_84 (.A(A[21]), .B(M_temp[21]), .ZN(n_63));
   XNOR2_X1 i_85 (.A(n_62), .B(n_63), .ZN(p_0[21]));
   INV_X1 i_86 (.A(A[21]), .ZN(n_64));
   AOI22_X1 i_87 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(M_temp[21]), .ZN(n_65));
   XOR2_X1 i_88 (.A(M_temp[22]), .B(A[22]), .Z(n_66));
   XNOR2_X1 i_89 (.A(n_65), .B(n_66), .ZN(p_0[22]));
   INV_X1 i_90 (.A(M_temp[22]), .ZN(n_67));
   OAI22_X1 i_91 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(A[22]), .ZN(n_68));
   XNOR2_X1 i_92 (.A(A[23]), .B(M_temp[23]), .ZN(n_69));
   XNOR2_X1 i_93 (.A(n_68), .B(n_69), .ZN(p_0[23]));
   INV_X1 i_94 (.A(A[23]), .ZN(n_70));
   AOI22_X1 i_95 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(M_temp[23]), .ZN(n_71));
   XOR2_X1 i_96 (.A(M_temp[24]), .B(A[24]), .Z(n_72));
   XNOR2_X1 i_97 (.A(n_71), .B(n_72), .ZN(p_0[24]));
   INV_X1 i_98 (.A(M_temp[24]), .ZN(n_73));
   OAI22_X1 i_99 (.A1(n_71), .A2(n_72), .B1(n_73), .B2(A[24]), .ZN(n_74));
   XNOR2_X1 i_100 (.A(A[25]), .B(M_temp[25]), .ZN(n_75));
   XNOR2_X1 i_101 (.A(n_74), .B(n_75), .ZN(p_0[25]));
   INV_X1 i_102 (.A(A[25]), .ZN(n_76));
   AOI22_X1 i_103 (.A1(n_74), .A2(n_75), .B1(n_76), .B2(M_temp[25]), .ZN(n_77));
   XOR2_X1 i_104 (.A(M_temp[26]), .B(A[26]), .Z(n_78));
   XNOR2_X1 i_105 (.A(n_77), .B(n_78), .ZN(p_0[26]));
   INV_X1 i_106 (.A(M_temp[26]), .ZN(n_79));
   OAI22_X1 i_107 (.A1(n_77), .A2(n_78), .B1(n_79), .B2(A[26]), .ZN(n_80));
   XNOR2_X1 i_108 (.A(A[27]), .B(M_temp[27]), .ZN(n_81));
   XNOR2_X1 i_109 (.A(n_80), .B(n_81), .ZN(p_0[27]));
   INV_X1 i_110 (.A(A[27]), .ZN(n_82));
   AOI22_X1 i_111 (.A1(n_80), .A2(n_81), .B1(n_82), .B2(M_temp[27]), .ZN(n_83));
   XOR2_X1 i_112 (.A(M_temp[28]), .B(A[28]), .Z(n_84));
   XNOR2_X1 i_113 (.A(n_83), .B(n_84), .ZN(p_0[28]));
   INV_X1 i_114 (.A(M_temp[28]), .ZN(n_85));
   OAI22_X1 i_115 (.A1(n_83), .A2(n_84), .B1(n_85), .B2(A[28]), .ZN(n_86));
   XNOR2_X1 i_116 (.A(A[29]), .B(M_temp[29]), .ZN(n_87));
   XNOR2_X1 i_117 (.A(n_86), .B(n_87), .ZN(p_0[29]));
   INV_X1 i_118 (.A(A[29]), .ZN(n_88));
   AOI22_X1 i_119 (.A1(n_86), .A2(n_87), .B1(n_88), .B2(M_temp[29]), .ZN(n_89));
   INV_X1 i_120 (.A(M_temp[30]), .ZN(n_90));
   OR2_X1 i_121 (.A1(n_90), .A2(A[30]), .ZN(n_91));
   NAND2_X1 i_122 (.A1(n_90), .A2(A[30]), .ZN(n_92));
   NAND2_X1 i_123 (.A1(n_91), .A2(n_92), .ZN(n_93));
   XNOR2_X1 i_124 (.A(n_89), .B(n_93), .ZN(p_0[30]));
   INV_X1 i_125 (.A(n_92), .ZN(n_94));
   AOI21_X1 i_126 (.A(n_94), .B1(n_89), .B2(n_91), .ZN(n_95));
   XNOR2_X1 i_127 (.A(A[31]), .B(M_temp[31]), .ZN(n_96));
   XNOR2_X1 i_128 (.A(n_95), .B(n_96), .ZN(p_0[31]));
endmodule

module datapath__0_0(M_temp, A, A0);
   input [31:0]M_temp;
   input [31:0]A;
   output [31:0]A0;

   HA_X1 i_0 (.A(M_temp[0]), .B(A[0]), .CO(n_0), .S(A0[0]));
   FA_X1 i_1 (.A(M_temp[1]), .B(A[1]), .CI(n_0), .CO(n_1), .S(A0[1]));
   FA_X1 i_2 (.A(M_temp[2]), .B(A[2]), .CI(n_1), .CO(n_2), .S(A0[2]));
   FA_X1 i_3 (.A(M_temp[3]), .B(A[3]), .CI(n_2), .CO(n_3), .S(A0[3]));
   FA_X1 i_4 (.A(M_temp[4]), .B(A[4]), .CI(n_3), .CO(n_4), .S(A0[4]));
   FA_X1 i_5 (.A(M_temp[5]), .B(A[5]), .CI(n_4), .CO(n_5), .S(A0[5]));
   FA_X1 i_6 (.A(M_temp[6]), .B(A[6]), .CI(n_5), .CO(n_6), .S(A0[6]));
   FA_X1 i_7 (.A(M_temp[7]), .B(A[7]), .CI(n_6), .CO(n_7), .S(A0[7]));
   FA_X1 i_8 (.A(M_temp[8]), .B(A[8]), .CI(n_7), .CO(n_8), .S(A0[8]));
   FA_X1 i_9 (.A(M_temp[9]), .B(A[9]), .CI(n_8), .CO(n_9), .S(A0[9]));
   FA_X1 i_10 (.A(M_temp[10]), .B(A[10]), .CI(n_9), .CO(n_10), .S(A0[10]));
   FA_X1 i_11 (.A(M_temp[11]), .B(A[11]), .CI(n_10), .CO(n_11), .S(A0[11]));
   FA_X1 i_12 (.A(M_temp[12]), .B(A[12]), .CI(n_11), .CO(n_12), .S(A0[12]));
   FA_X1 i_13 (.A(M_temp[13]), .B(A[13]), .CI(n_12), .CO(n_13), .S(A0[13]));
   FA_X1 i_14 (.A(M_temp[14]), .B(A[14]), .CI(n_13), .CO(n_14), .S(A0[14]));
   FA_X1 i_15 (.A(M_temp[15]), .B(A[15]), .CI(n_14), .CO(n_15), .S(A0[15]));
   FA_X1 i_16 (.A(M_temp[16]), .B(A[16]), .CI(n_15), .CO(n_16), .S(A0[16]));
   FA_X1 i_17 (.A(M_temp[17]), .B(A[17]), .CI(n_16), .CO(n_17), .S(A0[17]));
   FA_X1 i_18 (.A(M_temp[18]), .B(A[18]), .CI(n_17), .CO(n_18), .S(A0[18]));
   FA_X1 i_19 (.A(M_temp[19]), .B(A[19]), .CI(n_18), .CO(n_19), .S(A0[19]));
   FA_X1 i_20 (.A(M_temp[20]), .B(A[20]), .CI(n_19), .CO(n_20), .S(A0[20]));
   FA_X1 i_21 (.A(M_temp[21]), .B(A[21]), .CI(n_20), .CO(n_21), .S(A0[21]));
   FA_X1 i_22 (.A(M_temp[22]), .B(A[22]), .CI(n_21), .CO(n_22), .S(A0[22]));
   FA_X1 i_23 (.A(M_temp[23]), .B(A[23]), .CI(n_22), .CO(n_23), .S(A0[23]));
   FA_X1 i_24 (.A(M_temp[24]), .B(A[24]), .CI(n_23), .CO(n_24), .S(A0[24]));
   FA_X1 i_25 (.A(M_temp[25]), .B(A[25]), .CI(n_24), .CO(n_25), .S(A0[25]));
   FA_X1 i_26 (.A(M_temp[26]), .B(A[26]), .CI(n_25), .CO(n_26), .S(A0[26]));
   FA_X1 i_27 (.A(M_temp[27]), .B(A[27]), .CI(n_26), .CO(n_27), .S(A0[27]));
   FA_X1 i_28 (.A(M_temp[28]), .B(A[28]), .CI(n_27), .CO(n_28), .S(A0[28]));
   FA_X1 i_29 (.A(M_temp[29]), .B(A[29]), .CI(n_28), .CO(n_29), .S(A0[29]));
   FA_X1 i_30 (.A(M_temp[30]), .B(A[30]), .CI(n_29), .CO(n_30), .S(A0[30]));
   XNOR2_X1 i_31 (.A(M_temp[31]), .B(A[31]), .ZN(n_31));
   XNOR2_X1 i_32 (.A(n_31), .B(n_30), .ZN(A0[31]));
endmodule

module datapath__0_8(Count, p_0);
   input [31:0]Count;
   output [31:0]p_0;

   INV_X1 i_0 (.A(Count[0]), .ZN(p_0[0]));
   XNOR2_X1 i_1 (.A(Count[1]), .B(Count[0]), .ZN(p_0[1]));
   OR2_X1 i_2 (.A1(Count[1]), .A2(Count[0]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(Count[2]), .B(n_0), .ZN(p_0[2]));
   OR2_X1 i_4 (.A1(Count[2]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_5 (.A(Count[3]), .B(n_1), .ZN(p_0[3]));
   OR2_X1 i_6 (.A1(Count[3]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_7 (.A(Count[4]), .B(n_2), .ZN(p_0[4]));
   OR2_X1 i_8 (.A1(Count[4]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_9 (.A(Count[5]), .B(n_3), .ZN(p_0[5]));
   OR2_X1 i_10 (.A1(Count[5]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_11 (.A(Count[6]), .B(n_4), .ZN(p_0[6]));
   OR2_X1 i_12 (.A1(Count[6]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_13 (.A(Count[7]), .B(n_5), .ZN(p_0[7]));
   OR2_X1 i_14 (.A1(Count[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_15 (.A(Count[8]), .B(n_6), .ZN(p_0[8]));
   OR2_X1 i_16 (.A1(Count[8]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_17 (.A(Count[9]), .B(n_7), .ZN(p_0[9]));
   OR2_X1 i_18 (.A1(Count[9]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_19 (.A(Count[10]), .B(n_8), .ZN(p_0[10]));
   OR2_X1 i_20 (.A1(Count[10]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_21 (.A(Count[11]), .B(n_9), .ZN(p_0[11]));
   OR2_X1 i_22 (.A1(Count[11]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_23 (.A(Count[12]), .B(n_10), .ZN(p_0[12]));
   OR2_X1 i_24 (.A1(Count[12]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_25 (.A(Count[13]), .B(n_11), .ZN(p_0[13]));
   OR2_X1 i_26 (.A1(Count[13]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_27 (.A(Count[14]), .B(n_12), .ZN(p_0[14]));
   OR2_X1 i_28 (.A1(Count[14]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_29 (.A(Count[15]), .B(n_13), .ZN(p_0[15]));
   OR2_X1 i_30 (.A1(Count[15]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_31 (.A(Count[16]), .B(n_14), .ZN(p_0[16]));
   OR2_X1 i_32 (.A1(Count[16]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_33 (.A(Count[17]), .B(n_15), .ZN(p_0[17]));
   OR2_X1 i_34 (.A1(Count[17]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_35 (.A(Count[18]), .B(n_16), .ZN(p_0[18]));
   OR2_X1 i_36 (.A1(Count[18]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_37 (.A(Count[19]), .B(n_17), .ZN(p_0[19]));
   OR2_X1 i_38 (.A1(Count[19]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_39 (.A(Count[20]), .B(n_18), .ZN(p_0[20]));
   OR2_X1 i_40 (.A1(Count[20]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_41 (.A(Count[21]), .B(n_19), .ZN(p_0[21]));
   OR2_X1 i_42 (.A1(Count[21]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_43 (.A(Count[22]), .B(n_20), .ZN(p_0[22]));
   OR2_X1 i_44 (.A1(Count[22]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_45 (.A(Count[23]), .B(n_21), .ZN(p_0[23]));
   OR2_X1 i_46 (.A1(Count[23]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_47 (.A(Count[24]), .B(n_22), .ZN(p_0[24]));
   OR2_X1 i_48 (.A1(Count[24]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_49 (.A(Count[25]), .B(n_23), .ZN(p_0[25]));
   OR2_X1 i_50 (.A1(Count[25]), .A2(n_23), .ZN(n_24));
   XNOR2_X1 i_51 (.A(Count[26]), .B(n_24), .ZN(p_0[26]));
   OR2_X1 i_52 (.A1(Count[26]), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_53 (.A(Count[27]), .B(n_25), .ZN(p_0[27]));
   OR2_X1 i_54 (.A1(Count[27]), .A2(n_25), .ZN(n_26));
   XNOR2_X1 i_55 (.A(Count[28]), .B(n_26), .ZN(p_0[28]));
   OR2_X1 i_56 (.A1(Count[28]), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_57 (.A(Count[29]), .B(n_27), .ZN(p_0[29]));
   OR2_X1 i_58 (.A1(Count[29]), .A2(n_27), .ZN(n_28));
   XNOR2_X1 i_59 (.A(Count[30]), .B(n_28), .ZN(p_0[30]));
   OR2_X1 i_60 (.A1(Count[30]), .A2(n_28), .ZN(n_29));
   XNOR2_X1 i_61 (.A(Count[31]), .B(n_29), .ZN(p_0[31]));
endmodule

module both(clk, load, reset, M, Q, P);
   input clk;
   input load;
   input reset;
   input [31:0]M;
   input [31:0]Q;
   output [63:0]P;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_97;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_2_0;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_2_1;
   wire n_0_101;
   wire n_0_2_2;
   wire n_0_102;
   wire n_0_2_3;
   wire n_0_103;
   wire n_0_2_4;
   wire n_0_104;
   wire n_0_2_5;
   wire n_0_105;
   wire n_0_2_6;
   wire n_0_106;
   wire n_0_2_7;
   wire n_0_107;
   wire n_0_2_8;
   wire n_0_108;
   wire n_0_2_9;
   wire n_0_109;
   wire n_0_2_10;
   wire n_0_110;
   wire n_0_2_11;
   wire n_0_111;
   wire n_0_2_12;
   wire n_0_112;
   wire n_0_2_13;
   wire n_0_113;
   wire n_0_2_14;
   wire n_0_114;
   wire n_0_2_15;
   wire n_0_115;
   wire n_0_2_16;
   wire n_0_116;
   wire n_0_2_17;
   wire n_0_117;
   wire n_0_2_18;
   wire n_0_118;
   wire n_0_2_19;
   wire n_0_119;
   wire n_0_2_20;
   wire n_0_120;
   wire n_0_2_21;
   wire n_0_121;
   wire n_0_2_22;
   wire n_0_122;
   wire n_0_2_23;
   wire n_0_123;
   wire n_0_2_24;
   wire n_0_124;
   wire n_0_2_25;
   wire n_0_125;
   wire n_0_2_26;
   wire n_0_126;
   wire n_0_2_27;
   wire n_0_127;
   wire n_0_2_28;
   wire n_0_128;
   wire n_0_2_29;
   wire n_0_129;
   wire n_0_2_30;
   wire n_0_130;
   wire n_0_2_31;
   wire n_0_131;
   wire n_0_2_32;
   wire n_0_132;
   wire n_0_2_33;
   wire n_0_2_34;
   wire n_0_133;
   wire n_0_2_35;
   wire n_0_2_36;
   wire n_0_134;
   wire n_0_2_37;
   wire n_0_2_38;
   wire n_0_135;
   wire n_0_2_39;
   wire n_0_2_40;
   wire n_0_136;
   wire n_0_2_41;
   wire n_0_2_42;
   wire n_0_137;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_138;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_139;
   wire n_0_2_47;
   wire n_0_2_48;
   wire n_0_140;
   wire n_0_2_49;
   wire n_0_2_50;
   wire n_0_141;
   wire n_0_2_51;
   wire n_0_2_52;
   wire n_0_142;
   wire n_0_2_53;
   wire n_0_2_54;
   wire n_0_143;
   wire n_0_2_55;
   wire n_0_2_56;
   wire n_0_144;
   wire n_0_2_57;
   wire n_0_2_58;
   wire n_0_145;
   wire n_0_2_59;
   wire n_0_2_60;
   wire n_0_146;
   wire n_0_2_61;
   wire n_0_2_62;
   wire n_0_147;
   wire n_0_2_63;
   wire n_0_2_64;
   wire n_0_148;
   wire n_0_2_65;
   wire n_0_2_66;
   wire n_0_149;
   wire n_0_2_67;
   wire n_0_2_68;
   wire n_0_150;
   wire n_0_2_69;
   wire n_0_2_70;
   wire n_0_151;
   wire n_0_2_71;
   wire n_0_2_72;
   wire n_0_152;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_153;
   wire n_0_2_75;
   wire n_0_2_76;
   wire n_0_154;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_155;
   wire n_0_2_79;
   wire n_0_2_80;
   wire n_0_156;
   wire n_0_2_81;
   wire n_0_2_82;
   wire n_0_157;
   wire n_0_2_83;
   wire n_0_2_84;
   wire n_0_158;
   wire n_0_2_85;
   wire n_0_2_86;
   wire n_0_159;
   wire n_0_2_87;
   wire n_0_2_88;
   wire n_0_160;
   wire n_0_2_89;
   wire n_0_2_90;
   wire n_0_161;
   wire n_0_2_91;
   wire n_0_2_92;
   wire n_0_162;
   wire n_0_2_93;
   wire n_0_2_94;
   wire n_0_163;
   wire n_0_2_95;
   wire n_0_164;
   wire n_0_2_96;
   wire n_0_2_97;
   wire n_0_2_98;
   wire n_0_230;
   wire n_0_2_99;
   wire n_0_2_100;
   wire n_0_165;
   wire n_0_2_101;
   wire n_0_2_102;
   wire n_0_2_103;
   wire n_0_2_104;
   wire n_0_2_105;
   wire n_0_96;
   wire n_0_2_106;
   wire n_0_2_107;
   wire n_0_2_108;
   wire n_0_2_109;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_2_114;
   wire n_0_2_115;
   wire n_0_2_116;
   wire n_0_2_117;
   wire n_0_2_118;
   wire n_0_2_119;
   wire n_0_2_120;
   wire Q_minus_one;
   wire n_0_100;
   wire n_0_98;
   wire [31:0]Count;
   wire n_0_99;
   wire [31:0]M_temp;

   datapath i_0_0 (.A({P[63], P[62], P[61], P[60], P[59], P[58], P[57], P[56], 
      P[55], P[54], P[53], P[52], P[51], P[50], P[49], P[48], P[47], P[46], 
      P[45], P[44], P[43], P[42], P[41], P[40], P[39], P[38], P[37], P[36], 
      P[35], P[34], P[33], P[32]}), .p_0({n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, 
      n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}), .M_temp(
      M_temp));
   datapath__0_0 i_0_1 (.M_temp(M_temp), .A({P[63], P[62], P[61], P[60], P[59], 
      P[58], P[57], P[56], P[55], P[54], P[53], P[52], P[51], P[50], P[49], 
      P[48], P[47], P[46], P[45], P[44], P[43], P[42], P[41], P[40], P[39], 
      P[38], P[37], P[36], P[35], P[34], P[33], P[32]}), .A0({n_0_63, n_0_62, 
      n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, 
      n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, 
      n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
      n_0_34, n_0_33, n_0_32}));
   datapath__0_8 i_0_11 (.Count(Count), .p_0({n_0_197, n_0_196, n_0_195, n_0_194, 
      n_0_193, n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, 
      n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, 
      n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166}));
   AND2_X1 i_0_2_0 (.A1(n_0_2_118), .A2(M[0]), .ZN(n_0_64));
   AND2_X1 i_0_2_1 (.A1(n_0_2_118), .A2(M[1]), .ZN(n_0_65));
   AND2_X1 i_0_2_2 (.A1(n_0_2_118), .A2(M[2]), .ZN(n_0_66));
   AND2_X1 i_0_2_3 (.A1(n_0_2_118), .A2(M[3]), .ZN(n_0_67));
   AND2_X1 i_0_2_4 (.A1(n_0_2_118), .A2(M[4]), .ZN(n_0_68));
   AND2_X1 i_0_2_5 (.A1(n_0_2_118), .A2(M[5]), .ZN(n_0_69));
   AND2_X1 i_0_2_6 (.A1(n_0_2_118), .A2(M[6]), .ZN(n_0_70));
   AND2_X1 i_0_2_7 (.A1(n_0_2_118), .A2(M[7]), .ZN(n_0_71));
   AND2_X1 i_0_2_8 (.A1(n_0_2_118), .A2(M[8]), .ZN(n_0_72));
   AND2_X1 i_0_2_9 (.A1(n_0_2_118), .A2(M[9]), .ZN(n_0_73));
   AND2_X1 i_0_2_10 (.A1(n_0_2_118), .A2(M[10]), .ZN(n_0_74));
   AND2_X1 i_0_2_11 (.A1(n_0_2_118), .A2(M[11]), .ZN(n_0_75));
   AND2_X1 i_0_2_12 (.A1(n_0_2_118), .A2(M[12]), .ZN(n_0_76));
   AND2_X1 i_0_2_13 (.A1(n_0_2_118), .A2(M[13]), .ZN(n_0_77));
   AND2_X1 i_0_2_14 (.A1(n_0_2_118), .A2(M[14]), .ZN(n_0_78));
   AND2_X1 i_0_2_15 (.A1(n_0_2_118), .A2(M[15]), .ZN(n_0_79));
   AND2_X1 i_0_2_16 (.A1(n_0_2_118), .A2(M[16]), .ZN(n_0_80));
   AND2_X1 i_0_2_17 (.A1(n_0_2_118), .A2(M[17]), .ZN(n_0_81));
   AND2_X1 i_0_2_18 (.A1(n_0_2_118), .A2(M[18]), .ZN(n_0_82));
   AND2_X1 i_0_2_19 (.A1(n_0_2_118), .A2(M[19]), .ZN(n_0_83));
   AND2_X1 i_0_2_20 (.A1(n_0_2_118), .A2(M[20]), .ZN(n_0_84));
   AND2_X1 i_0_2_21 (.A1(n_0_2_118), .A2(M[21]), .ZN(n_0_85));
   AND2_X1 i_0_2_22 (.A1(n_0_2_118), .A2(M[22]), .ZN(n_0_86));
   AND2_X1 i_0_2_23 (.A1(n_0_2_118), .A2(M[23]), .ZN(n_0_87));
   AND2_X1 i_0_2_24 (.A1(n_0_2_118), .A2(M[24]), .ZN(n_0_88));
   AND2_X1 i_0_2_25 (.A1(n_0_2_118), .A2(M[25]), .ZN(n_0_89));
   AND2_X1 i_0_2_26 (.A1(n_0_2_118), .A2(M[26]), .ZN(n_0_90));
   AND2_X1 i_0_2_27 (.A1(n_0_2_118), .A2(M[27]), .ZN(n_0_91));
   AND2_X1 i_0_2_28 (.A1(n_0_2_118), .A2(M[28]), .ZN(n_0_92));
   AND2_X1 i_0_2_29 (.A1(n_0_2_118), .A2(M[29]), .ZN(n_0_93));
   AND2_X1 i_0_2_30 (.A1(n_0_2_118), .A2(M[30]), .ZN(n_0_94));
   AND2_X1 i_0_2_31 (.A1(n_0_2_118), .A2(M[31]), .ZN(n_0_95));
   NOR2_X1 i_0_2_32 (.A1(n_0_2_119), .A2(reset), .ZN(n_0_97));
   AND2_X1 i_0_2_33 (.A1(n_0_166), .A2(n_0_2_1), .ZN(n_0_198));
   AND2_X1 i_0_2_34 (.A1(n_0_167), .A2(n_0_2_1), .ZN(n_0_199));
   AND2_X1 i_0_2_35 (.A1(n_0_168), .A2(n_0_2_1), .ZN(n_0_200));
   AND2_X1 i_0_2_36 (.A1(n_0_169), .A2(n_0_2_1), .ZN(n_0_201));
   AND2_X1 i_0_2_37 (.A1(n_0_170), .A2(n_0_2_1), .ZN(n_0_202));
   INV_X1 i_0_2_38 (.A(n_0_2_0), .ZN(n_0_203));
   AOI21_X1 i_0_2_39 (.A(reset), .B1(n_0_171), .B2(n_0_2_106), .ZN(n_0_2_0));
   AND2_X1 i_0_2_40 (.A1(n_0_172), .A2(n_0_2_1), .ZN(n_0_204));
   AND2_X1 i_0_2_41 (.A1(n_0_173), .A2(n_0_2_1), .ZN(n_0_205));
   AND2_X1 i_0_2_42 (.A1(n_0_174), .A2(n_0_2_1), .ZN(n_0_206));
   AND2_X1 i_0_2_43 (.A1(n_0_175), .A2(n_0_2_1), .ZN(n_0_207));
   AND2_X1 i_0_2_44 (.A1(n_0_176), .A2(n_0_2_1), .ZN(n_0_208));
   AND2_X1 i_0_2_45 (.A1(n_0_177), .A2(n_0_2_1), .ZN(n_0_209));
   AND2_X1 i_0_2_46 (.A1(n_0_178), .A2(n_0_2_1), .ZN(n_0_210));
   AND2_X1 i_0_2_47 (.A1(n_0_179), .A2(n_0_2_1), .ZN(n_0_211));
   AND2_X1 i_0_2_48 (.A1(n_0_180), .A2(n_0_2_1), .ZN(n_0_212));
   AND2_X1 i_0_2_49 (.A1(n_0_181), .A2(n_0_2_1), .ZN(n_0_213));
   AND2_X1 i_0_2_50 (.A1(n_0_182), .A2(n_0_2_1), .ZN(n_0_214));
   AND2_X1 i_0_2_51 (.A1(n_0_183), .A2(n_0_2_1), .ZN(n_0_215));
   AND2_X1 i_0_2_52 (.A1(n_0_184), .A2(n_0_2_1), .ZN(n_0_216));
   AND2_X1 i_0_2_53 (.A1(n_0_185), .A2(n_0_2_1), .ZN(n_0_217));
   AND2_X1 i_0_2_54 (.A1(n_0_186), .A2(n_0_2_1), .ZN(n_0_218));
   AND2_X1 i_0_2_55 (.A1(n_0_187), .A2(n_0_2_1), .ZN(n_0_219));
   AND2_X1 i_0_2_56 (.A1(n_0_188), .A2(n_0_2_1), .ZN(n_0_220));
   AND2_X1 i_0_2_57 (.A1(n_0_189), .A2(n_0_2_1), .ZN(n_0_221));
   AND2_X1 i_0_2_58 (.A1(n_0_190), .A2(n_0_2_1), .ZN(n_0_222));
   AND2_X1 i_0_2_59 (.A1(n_0_191), .A2(n_0_2_1), .ZN(n_0_223));
   AND2_X1 i_0_2_60 (.A1(n_0_192), .A2(n_0_2_1), .ZN(n_0_224));
   AND2_X1 i_0_2_61 (.A1(n_0_193), .A2(n_0_2_1), .ZN(n_0_225));
   AND2_X1 i_0_2_62 (.A1(n_0_194), .A2(n_0_2_1), .ZN(n_0_226));
   AND2_X1 i_0_2_63 (.A1(n_0_195), .A2(n_0_2_1), .ZN(n_0_227));
   AND2_X1 i_0_2_64 (.A1(n_0_196), .A2(n_0_2_1), .ZN(n_0_228));
   AND2_X1 i_0_2_65 (.A1(n_0_197), .A2(n_0_2_1), .ZN(n_0_229));
   NOR2_X1 i_0_2_66 (.A1(reset), .A2(n_0_2_107), .ZN(n_0_2_1));
   INV_X1 i_0_2_67 (.A(n_0_2_2), .ZN(n_0_101));
   AOI222_X1 i_0_2_68 (.A1(Q[0]), .A2(n_0_2_100), .B1(P[1]), .B2(n_0_2_105), 
      .C1(P[0]), .C2(n_0_2_99), .ZN(n_0_2_2));
   INV_X1 i_0_2_69 (.A(n_0_2_3), .ZN(n_0_102));
   AOI222_X1 i_0_2_70 (.A1(Q[1]), .A2(n_0_2_100), .B1(P[2]), .B2(n_0_2_105), 
      .C1(P[1]), .C2(n_0_2_99), .ZN(n_0_2_3));
   INV_X1 i_0_2_71 (.A(n_0_2_4), .ZN(n_0_103));
   AOI222_X1 i_0_2_72 (.A1(Q[2]), .A2(n_0_2_100), .B1(P[3]), .B2(n_0_2_105), 
      .C1(P[2]), .C2(n_0_2_99), .ZN(n_0_2_4));
   INV_X1 i_0_2_73 (.A(n_0_2_5), .ZN(n_0_104));
   AOI222_X1 i_0_2_74 (.A1(Q[3]), .A2(n_0_2_100), .B1(P[4]), .B2(n_0_2_105), 
      .C1(P[3]), .C2(n_0_2_99), .ZN(n_0_2_5));
   INV_X1 i_0_2_75 (.A(n_0_2_6), .ZN(n_0_105));
   AOI222_X1 i_0_2_76 (.A1(Q[4]), .A2(n_0_2_100), .B1(P[5]), .B2(n_0_2_105), 
      .C1(P[4]), .C2(n_0_2_99), .ZN(n_0_2_6));
   INV_X1 i_0_2_77 (.A(n_0_2_7), .ZN(n_0_106));
   AOI222_X1 i_0_2_78 (.A1(Q[5]), .A2(n_0_2_100), .B1(P[6]), .B2(n_0_2_105), 
      .C1(P[5]), .C2(n_0_2_99), .ZN(n_0_2_7));
   INV_X1 i_0_2_79 (.A(n_0_2_8), .ZN(n_0_107));
   AOI222_X1 i_0_2_80 (.A1(Q[6]), .A2(n_0_2_100), .B1(P[7]), .B2(n_0_2_105), 
      .C1(P[6]), .C2(n_0_2_99), .ZN(n_0_2_8));
   INV_X1 i_0_2_81 (.A(n_0_2_9), .ZN(n_0_108));
   AOI222_X1 i_0_2_82 (.A1(Q[7]), .A2(n_0_2_100), .B1(P[8]), .B2(n_0_2_105), 
      .C1(P[7]), .C2(n_0_2_99), .ZN(n_0_2_9));
   INV_X1 i_0_2_83 (.A(n_0_2_10), .ZN(n_0_109));
   AOI222_X1 i_0_2_84 (.A1(Q[8]), .A2(n_0_2_100), .B1(P[9]), .B2(n_0_2_105), 
      .C1(P[8]), .C2(n_0_2_99), .ZN(n_0_2_10));
   INV_X1 i_0_2_85 (.A(n_0_2_11), .ZN(n_0_110));
   AOI222_X1 i_0_2_86 (.A1(Q[9]), .A2(n_0_2_100), .B1(P[10]), .B2(n_0_2_105), 
      .C1(P[9]), .C2(n_0_2_99), .ZN(n_0_2_11));
   INV_X1 i_0_2_87 (.A(n_0_2_12), .ZN(n_0_111));
   AOI222_X1 i_0_2_88 (.A1(Q[10]), .A2(n_0_2_100), .B1(P[11]), .B2(n_0_2_105), 
      .C1(P[10]), .C2(n_0_2_99), .ZN(n_0_2_12));
   INV_X1 i_0_2_89 (.A(n_0_2_13), .ZN(n_0_112));
   AOI222_X1 i_0_2_90 (.A1(Q[11]), .A2(n_0_2_100), .B1(P[12]), .B2(n_0_2_105), 
      .C1(P[11]), .C2(n_0_2_99), .ZN(n_0_2_13));
   INV_X1 i_0_2_91 (.A(n_0_2_14), .ZN(n_0_113));
   AOI222_X1 i_0_2_92 (.A1(Q[12]), .A2(n_0_2_100), .B1(P[13]), .B2(n_0_2_105), 
      .C1(P[12]), .C2(n_0_2_99), .ZN(n_0_2_14));
   INV_X1 i_0_2_93 (.A(n_0_2_15), .ZN(n_0_114));
   AOI222_X1 i_0_2_94 (.A1(Q[13]), .A2(n_0_2_100), .B1(P[14]), .B2(n_0_2_105), 
      .C1(P[13]), .C2(n_0_2_99), .ZN(n_0_2_15));
   INV_X1 i_0_2_95 (.A(n_0_2_16), .ZN(n_0_115));
   AOI222_X1 i_0_2_96 (.A1(Q[14]), .A2(n_0_2_100), .B1(P[15]), .B2(n_0_2_105), 
      .C1(P[14]), .C2(n_0_2_99), .ZN(n_0_2_16));
   INV_X1 i_0_2_97 (.A(n_0_2_17), .ZN(n_0_116));
   AOI222_X1 i_0_2_98 (.A1(Q[15]), .A2(n_0_2_100), .B1(P[16]), .B2(n_0_2_105), 
      .C1(P[15]), .C2(n_0_2_99), .ZN(n_0_2_17));
   INV_X1 i_0_2_99 (.A(n_0_2_18), .ZN(n_0_117));
   AOI222_X1 i_0_2_100 (.A1(Q[16]), .A2(n_0_2_100), .B1(P[17]), .B2(n_0_2_105), 
      .C1(P[16]), .C2(n_0_2_99), .ZN(n_0_2_18));
   INV_X1 i_0_2_101 (.A(n_0_2_19), .ZN(n_0_118));
   AOI222_X1 i_0_2_102 (.A1(Q[17]), .A2(n_0_2_100), .B1(P[18]), .B2(n_0_2_105), 
      .C1(P[17]), .C2(n_0_2_99), .ZN(n_0_2_19));
   INV_X1 i_0_2_103 (.A(n_0_2_20), .ZN(n_0_119));
   AOI222_X1 i_0_2_104 (.A1(Q[18]), .A2(n_0_2_100), .B1(P[19]), .B2(n_0_2_105), 
      .C1(P[18]), .C2(n_0_2_99), .ZN(n_0_2_20));
   INV_X1 i_0_2_105 (.A(n_0_2_21), .ZN(n_0_120));
   AOI222_X1 i_0_2_106 (.A1(Q[19]), .A2(n_0_2_100), .B1(P[20]), .B2(n_0_2_105), 
      .C1(P[19]), .C2(n_0_2_99), .ZN(n_0_2_21));
   INV_X1 i_0_2_107 (.A(n_0_2_22), .ZN(n_0_121));
   AOI222_X1 i_0_2_108 (.A1(Q[20]), .A2(n_0_2_100), .B1(P[21]), .B2(n_0_2_105), 
      .C1(P[20]), .C2(n_0_2_99), .ZN(n_0_2_22));
   INV_X1 i_0_2_109 (.A(n_0_2_23), .ZN(n_0_122));
   AOI222_X1 i_0_2_110 (.A1(Q[21]), .A2(n_0_2_100), .B1(P[22]), .B2(n_0_2_105), 
      .C1(P[21]), .C2(n_0_2_99), .ZN(n_0_2_23));
   INV_X1 i_0_2_111 (.A(n_0_2_24), .ZN(n_0_123));
   AOI222_X1 i_0_2_112 (.A1(Q[22]), .A2(n_0_2_100), .B1(P[23]), .B2(n_0_2_105), 
      .C1(P[22]), .C2(n_0_2_99), .ZN(n_0_2_24));
   INV_X1 i_0_2_113 (.A(n_0_2_25), .ZN(n_0_124));
   AOI222_X1 i_0_2_114 (.A1(Q[23]), .A2(n_0_2_100), .B1(P[24]), .B2(n_0_2_105), 
      .C1(P[23]), .C2(n_0_2_99), .ZN(n_0_2_25));
   INV_X1 i_0_2_115 (.A(n_0_2_26), .ZN(n_0_125));
   AOI222_X1 i_0_2_116 (.A1(Q[24]), .A2(n_0_2_100), .B1(P[25]), .B2(n_0_2_105), 
      .C1(P[24]), .C2(n_0_2_99), .ZN(n_0_2_26));
   INV_X1 i_0_2_117 (.A(n_0_2_27), .ZN(n_0_126));
   AOI222_X1 i_0_2_118 (.A1(Q[25]), .A2(n_0_2_100), .B1(P[26]), .B2(n_0_2_105), 
      .C1(P[25]), .C2(n_0_2_99), .ZN(n_0_2_27));
   INV_X1 i_0_2_119 (.A(n_0_2_28), .ZN(n_0_127));
   AOI222_X1 i_0_2_120 (.A1(Q[26]), .A2(n_0_2_100), .B1(P[27]), .B2(n_0_2_105), 
      .C1(P[26]), .C2(n_0_2_99), .ZN(n_0_2_28));
   INV_X1 i_0_2_121 (.A(n_0_2_29), .ZN(n_0_128));
   AOI222_X1 i_0_2_122 (.A1(Q[27]), .A2(n_0_2_100), .B1(P[28]), .B2(n_0_2_105), 
      .C1(P[27]), .C2(n_0_2_99), .ZN(n_0_2_29));
   INV_X1 i_0_2_123 (.A(n_0_2_30), .ZN(n_0_129));
   AOI222_X1 i_0_2_124 (.A1(Q[28]), .A2(n_0_2_100), .B1(P[29]), .B2(n_0_2_105), 
      .C1(P[28]), .C2(n_0_2_99), .ZN(n_0_2_30));
   INV_X1 i_0_2_125 (.A(n_0_2_31), .ZN(n_0_130));
   AOI222_X1 i_0_2_126 (.A1(Q[29]), .A2(n_0_2_100), .B1(P[30]), .B2(n_0_2_105), 
      .C1(P[29]), .C2(n_0_2_99), .ZN(n_0_2_31));
   INV_X1 i_0_2_127 (.A(n_0_2_32), .ZN(n_0_131));
   AOI222_X1 i_0_2_128 (.A1(Q[30]), .A2(n_0_2_100), .B1(P[31]), .B2(n_0_2_105), 
      .C1(P[30]), .C2(n_0_2_99), .ZN(n_0_2_32));
   NAND2_X1 i_0_2_129 (.A1(n_0_2_34), .A2(n_0_2_33), .ZN(n_0_132));
   AOI22_X1 i_0_2_130 (.A1(n_0_0), .A2(n_0_2_102), .B1(P[32]), .B2(n_0_2_97), 
      .ZN(n_0_2_33));
   AOI222_X1 i_0_2_131 (.A1(P[31]), .A2(n_0_2_99), .B1(Q[31]), .B2(n_0_2_100), 
      .C1(n_0_32), .C2(n_0_2_103), .ZN(n_0_2_34));
   NAND2_X1 i_0_2_132 (.A1(n_0_2_36), .A2(n_0_2_35), .ZN(n_0_133));
   AOI22_X1 i_0_2_133 (.A1(n_0_1), .A2(n_0_2_102), .B1(P[32]), .B2(n_0_2_98), 
      .ZN(n_0_2_35));
   AOI22_X1 i_0_2_134 (.A1(n_0_33), .A2(n_0_2_103), .B1(P[33]), .B2(n_0_2_97), 
      .ZN(n_0_2_36));
   NAND2_X1 i_0_2_135 (.A1(n_0_2_38), .A2(n_0_2_37), .ZN(n_0_134));
   AOI22_X1 i_0_2_136 (.A1(n_0_2), .A2(n_0_2_102), .B1(P[33]), .B2(n_0_2_98), 
      .ZN(n_0_2_37));
   AOI22_X1 i_0_2_137 (.A1(n_0_34), .A2(n_0_2_103), .B1(P[34]), .B2(n_0_2_97), 
      .ZN(n_0_2_38));
   NAND2_X1 i_0_2_138 (.A1(n_0_2_40), .A2(n_0_2_39), .ZN(n_0_135));
   AOI22_X1 i_0_2_139 (.A1(n_0_3), .A2(n_0_2_102), .B1(P[34]), .B2(n_0_2_98), 
      .ZN(n_0_2_39));
   AOI22_X1 i_0_2_140 (.A1(n_0_35), .A2(n_0_2_103), .B1(P[35]), .B2(n_0_2_97), 
      .ZN(n_0_2_40));
   NAND2_X1 i_0_2_141 (.A1(n_0_2_42), .A2(n_0_2_41), .ZN(n_0_136));
   AOI22_X1 i_0_2_142 (.A1(n_0_4), .A2(n_0_2_102), .B1(P[35]), .B2(n_0_2_98), 
      .ZN(n_0_2_41));
   AOI22_X1 i_0_2_143 (.A1(n_0_36), .A2(n_0_2_103), .B1(P[36]), .B2(n_0_2_97), 
      .ZN(n_0_2_42));
   NAND2_X1 i_0_2_144 (.A1(n_0_2_44), .A2(n_0_2_43), .ZN(n_0_137));
   AOI22_X1 i_0_2_145 (.A1(n_0_5), .A2(n_0_2_102), .B1(P[36]), .B2(n_0_2_98), 
      .ZN(n_0_2_43));
   AOI22_X1 i_0_2_146 (.A1(n_0_37), .A2(n_0_2_103), .B1(P[37]), .B2(n_0_2_97), 
      .ZN(n_0_2_44));
   NAND2_X1 i_0_2_147 (.A1(n_0_2_46), .A2(n_0_2_45), .ZN(n_0_138));
   AOI22_X1 i_0_2_148 (.A1(n_0_6), .A2(n_0_2_102), .B1(P[37]), .B2(n_0_2_98), 
      .ZN(n_0_2_45));
   AOI22_X1 i_0_2_149 (.A1(n_0_38), .A2(n_0_2_103), .B1(P[38]), .B2(n_0_2_97), 
      .ZN(n_0_2_46));
   NAND2_X1 i_0_2_150 (.A1(n_0_2_48), .A2(n_0_2_47), .ZN(n_0_139));
   AOI22_X1 i_0_2_151 (.A1(n_0_7), .A2(n_0_2_102), .B1(P[38]), .B2(n_0_2_98), 
      .ZN(n_0_2_47));
   AOI22_X1 i_0_2_152 (.A1(n_0_39), .A2(n_0_2_103), .B1(P[39]), .B2(n_0_2_97), 
      .ZN(n_0_2_48));
   NAND2_X1 i_0_2_153 (.A1(n_0_2_50), .A2(n_0_2_49), .ZN(n_0_140));
   AOI22_X1 i_0_2_154 (.A1(n_0_8), .A2(n_0_2_102), .B1(P[39]), .B2(n_0_2_98), 
      .ZN(n_0_2_49));
   AOI22_X1 i_0_2_155 (.A1(n_0_40), .A2(n_0_2_103), .B1(P[40]), .B2(n_0_2_97), 
      .ZN(n_0_2_50));
   NAND2_X1 i_0_2_156 (.A1(n_0_2_52), .A2(n_0_2_51), .ZN(n_0_141));
   AOI22_X1 i_0_2_157 (.A1(n_0_9), .A2(n_0_2_102), .B1(P[40]), .B2(n_0_2_98), 
      .ZN(n_0_2_51));
   AOI22_X1 i_0_2_158 (.A1(n_0_41), .A2(n_0_2_103), .B1(P[41]), .B2(n_0_2_97), 
      .ZN(n_0_2_52));
   NAND2_X1 i_0_2_159 (.A1(n_0_2_54), .A2(n_0_2_53), .ZN(n_0_142));
   AOI22_X1 i_0_2_160 (.A1(n_0_10), .A2(n_0_2_102), .B1(P[41]), .B2(n_0_2_98), 
      .ZN(n_0_2_53));
   AOI22_X1 i_0_2_161 (.A1(n_0_42), .A2(n_0_2_103), .B1(P[42]), .B2(n_0_2_97), 
      .ZN(n_0_2_54));
   NAND2_X1 i_0_2_162 (.A1(n_0_2_56), .A2(n_0_2_55), .ZN(n_0_143));
   AOI22_X1 i_0_2_163 (.A1(n_0_11), .A2(n_0_2_102), .B1(P[42]), .B2(n_0_2_98), 
      .ZN(n_0_2_55));
   AOI22_X1 i_0_2_164 (.A1(n_0_43), .A2(n_0_2_103), .B1(P[43]), .B2(n_0_2_97), 
      .ZN(n_0_2_56));
   NAND2_X1 i_0_2_165 (.A1(n_0_2_58), .A2(n_0_2_57), .ZN(n_0_144));
   AOI22_X1 i_0_2_166 (.A1(n_0_12), .A2(n_0_2_102), .B1(P[43]), .B2(n_0_2_98), 
      .ZN(n_0_2_57));
   AOI22_X1 i_0_2_167 (.A1(n_0_44), .A2(n_0_2_103), .B1(P[44]), .B2(n_0_2_97), 
      .ZN(n_0_2_58));
   NAND2_X1 i_0_2_168 (.A1(n_0_2_60), .A2(n_0_2_59), .ZN(n_0_145));
   AOI22_X1 i_0_2_169 (.A1(n_0_13), .A2(n_0_2_102), .B1(P[44]), .B2(n_0_2_98), 
      .ZN(n_0_2_59));
   AOI22_X1 i_0_2_170 (.A1(n_0_45), .A2(n_0_2_103), .B1(P[45]), .B2(n_0_2_97), 
      .ZN(n_0_2_60));
   NAND2_X1 i_0_2_171 (.A1(n_0_2_62), .A2(n_0_2_61), .ZN(n_0_146));
   AOI22_X1 i_0_2_172 (.A1(n_0_14), .A2(n_0_2_102), .B1(P[45]), .B2(n_0_2_98), 
      .ZN(n_0_2_61));
   AOI22_X1 i_0_2_173 (.A1(n_0_46), .A2(n_0_2_103), .B1(P[46]), .B2(n_0_2_97), 
      .ZN(n_0_2_62));
   NAND2_X1 i_0_2_174 (.A1(n_0_2_64), .A2(n_0_2_63), .ZN(n_0_147));
   AOI22_X1 i_0_2_175 (.A1(n_0_15), .A2(n_0_2_102), .B1(P[46]), .B2(n_0_2_98), 
      .ZN(n_0_2_63));
   AOI22_X1 i_0_2_176 (.A1(n_0_47), .A2(n_0_2_103), .B1(P[47]), .B2(n_0_2_97), 
      .ZN(n_0_2_64));
   NAND2_X1 i_0_2_177 (.A1(n_0_2_66), .A2(n_0_2_65), .ZN(n_0_148));
   AOI22_X1 i_0_2_178 (.A1(P[47]), .A2(n_0_2_98), .B1(P[48]), .B2(n_0_2_97), 
      .ZN(n_0_2_65));
   AOI22_X1 i_0_2_179 (.A1(n_0_48), .A2(n_0_2_103), .B1(n_0_16), .B2(n_0_2_102), 
      .ZN(n_0_2_66));
   NAND2_X1 i_0_2_180 (.A1(n_0_2_68), .A2(n_0_2_67), .ZN(n_0_149));
   AOI22_X1 i_0_2_181 (.A1(P[48]), .A2(n_0_2_98), .B1(P[49]), .B2(n_0_2_97), 
      .ZN(n_0_2_67));
   AOI22_X1 i_0_2_182 (.A1(n_0_49), .A2(n_0_2_103), .B1(n_0_17), .B2(n_0_2_102), 
      .ZN(n_0_2_68));
   NAND2_X1 i_0_2_183 (.A1(n_0_2_70), .A2(n_0_2_69), .ZN(n_0_150));
   AOI22_X1 i_0_2_184 (.A1(n_0_18), .A2(n_0_2_102), .B1(P[49]), .B2(n_0_2_98), 
      .ZN(n_0_2_69));
   AOI22_X1 i_0_2_185 (.A1(n_0_50), .A2(n_0_2_103), .B1(P[50]), .B2(n_0_2_97), 
      .ZN(n_0_2_70));
   NAND2_X1 i_0_2_186 (.A1(n_0_2_72), .A2(n_0_2_71), .ZN(n_0_151));
   AOI22_X1 i_0_2_187 (.A1(n_0_19), .A2(n_0_2_102), .B1(P[50]), .B2(n_0_2_98), 
      .ZN(n_0_2_71));
   AOI22_X1 i_0_2_188 (.A1(n_0_51), .A2(n_0_2_103), .B1(P[51]), .B2(n_0_2_97), 
      .ZN(n_0_2_72));
   NAND2_X1 i_0_2_189 (.A1(n_0_2_74), .A2(n_0_2_73), .ZN(n_0_152));
   AOI22_X1 i_0_2_190 (.A1(n_0_20), .A2(n_0_2_102), .B1(P[51]), .B2(n_0_2_98), 
      .ZN(n_0_2_73));
   AOI22_X1 i_0_2_191 (.A1(n_0_52), .A2(n_0_2_103), .B1(P[52]), .B2(n_0_2_97), 
      .ZN(n_0_2_74));
   NAND2_X1 i_0_2_192 (.A1(n_0_2_76), .A2(n_0_2_75), .ZN(n_0_153));
   AOI22_X1 i_0_2_193 (.A1(n_0_21), .A2(n_0_2_102), .B1(P[52]), .B2(n_0_2_98), 
      .ZN(n_0_2_75));
   AOI22_X1 i_0_2_194 (.A1(n_0_53), .A2(n_0_2_103), .B1(P[53]), .B2(n_0_2_97), 
      .ZN(n_0_2_76));
   NAND2_X1 i_0_2_195 (.A1(n_0_2_78), .A2(n_0_2_77), .ZN(n_0_154));
   AOI22_X1 i_0_2_196 (.A1(n_0_22), .A2(n_0_2_102), .B1(P[53]), .B2(n_0_2_98), 
      .ZN(n_0_2_77));
   AOI22_X1 i_0_2_197 (.A1(n_0_54), .A2(n_0_2_103), .B1(P[54]), .B2(n_0_2_97), 
      .ZN(n_0_2_78));
   NAND2_X1 i_0_2_198 (.A1(n_0_2_80), .A2(n_0_2_79), .ZN(n_0_155));
   AOI22_X1 i_0_2_199 (.A1(n_0_23), .A2(n_0_2_102), .B1(P[54]), .B2(n_0_2_98), 
      .ZN(n_0_2_79));
   AOI22_X1 i_0_2_200 (.A1(n_0_55), .A2(n_0_2_103), .B1(P[55]), .B2(n_0_2_97), 
      .ZN(n_0_2_80));
   NAND2_X1 i_0_2_201 (.A1(n_0_2_82), .A2(n_0_2_81), .ZN(n_0_156));
   AOI22_X1 i_0_2_202 (.A1(n_0_24), .A2(n_0_2_102), .B1(P[55]), .B2(n_0_2_98), 
      .ZN(n_0_2_81));
   AOI22_X1 i_0_2_203 (.A1(n_0_56), .A2(n_0_2_103), .B1(P[56]), .B2(n_0_2_97), 
      .ZN(n_0_2_82));
   NAND2_X1 i_0_2_204 (.A1(n_0_2_84), .A2(n_0_2_83), .ZN(n_0_157));
   AOI22_X1 i_0_2_205 (.A1(n_0_25), .A2(n_0_2_102), .B1(P[56]), .B2(n_0_2_98), 
      .ZN(n_0_2_83));
   AOI22_X1 i_0_2_206 (.A1(n_0_57), .A2(n_0_2_103), .B1(P[57]), .B2(n_0_2_97), 
      .ZN(n_0_2_84));
   NAND2_X1 i_0_2_207 (.A1(n_0_2_86), .A2(n_0_2_85), .ZN(n_0_158));
   AOI22_X1 i_0_2_208 (.A1(n_0_26), .A2(n_0_2_102), .B1(P[57]), .B2(n_0_2_98), 
      .ZN(n_0_2_85));
   AOI22_X1 i_0_2_209 (.A1(n_0_58), .A2(n_0_2_103), .B1(P[58]), .B2(n_0_2_97), 
      .ZN(n_0_2_86));
   NAND2_X1 i_0_2_210 (.A1(n_0_2_88), .A2(n_0_2_87), .ZN(n_0_159));
   AOI22_X1 i_0_2_211 (.A1(n_0_27), .A2(n_0_2_102), .B1(P[58]), .B2(n_0_2_98), 
      .ZN(n_0_2_87));
   AOI22_X1 i_0_2_212 (.A1(n_0_59), .A2(n_0_2_103), .B1(P[59]), .B2(n_0_2_97), 
      .ZN(n_0_2_88));
   NAND2_X1 i_0_2_213 (.A1(n_0_2_90), .A2(n_0_2_89), .ZN(n_0_160));
   AOI22_X1 i_0_2_214 (.A1(n_0_28), .A2(n_0_2_102), .B1(P[59]), .B2(n_0_2_98), 
      .ZN(n_0_2_89));
   AOI22_X1 i_0_2_215 (.A1(n_0_60), .A2(n_0_2_103), .B1(P[60]), .B2(n_0_2_97), 
      .ZN(n_0_2_90));
   NAND2_X1 i_0_2_216 (.A1(n_0_2_92), .A2(n_0_2_91), .ZN(n_0_161));
   AOI22_X1 i_0_2_217 (.A1(n_0_29), .A2(n_0_2_102), .B1(P[60]), .B2(n_0_2_98), 
      .ZN(n_0_2_91));
   AOI22_X1 i_0_2_218 (.A1(n_0_61), .A2(n_0_2_103), .B1(P[61]), .B2(n_0_2_97), 
      .ZN(n_0_2_92));
   NAND2_X1 i_0_2_219 (.A1(n_0_2_94), .A2(n_0_2_93), .ZN(n_0_162));
   AOI22_X1 i_0_2_220 (.A1(n_0_30), .A2(n_0_2_102), .B1(P[61]), .B2(n_0_2_98), 
      .ZN(n_0_2_93));
   AOI22_X1 i_0_2_221 (.A1(n_0_62), .A2(n_0_2_103), .B1(P[62]), .B2(n_0_2_97), 
      .ZN(n_0_2_94));
   NAND2_X1 i_0_2_222 (.A1(n_0_2_101), .A2(n_0_2_95), .ZN(n_0_163));
   AOI22_X1 i_0_2_223 (.A1(P[62]), .A2(n_0_2_98), .B1(P[63]), .B2(n_0_2_97), 
      .ZN(n_0_2_95));
   NAND2_X1 i_0_2_224 (.A1(n_0_2_101), .A2(n_0_2_96), .ZN(n_0_164));
   OAI21_X1 i_0_2_225 (.A(P[63]), .B1(n_0_2_98), .B2(n_0_2_97), .ZN(n_0_2_96));
   AOI221_X1 i_0_2_226 (.A(n_0_2_104), .B1(Q_minus_one), .B2(n_0_2_119), 
      .C1(n_0_2_120), .C2(P[0]), .ZN(n_0_2_97));
   INV_X1 i_0_2_227 (.A(n_0_230), .ZN(n_0_2_98));
   NOR2_X1 i_0_2_228 (.A1(n_0_2_100), .A2(n_0_2_99), .ZN(n_0_230));
   NOR2_X1 i_0_2_229 (.A1(n_0_2_106), .A2(n_0_96), .ZN(n_0_2_99));
   INV_X1 i_0_2_230 (.A(n_0_165), .ZN(n_0_2_100));
   NAND2_X1 i_0_2_231 (.A1(n_0_2_118), .A2(load), .ZN(n_0_165));
   AOI22_X1 i_0_2_232 (.A1(n_0_63), .A2(n_0_2_103), .B1(n_0_31), .B2(n_0_2_102), 
      .ZN(n_0_2_101));
   NOR3_X1 i_0_2_233 (.A1(Q_minus_one), .A2(n_0_2_119), .A3(n_0_2_104), .ZN(
      n_0_2_102));
   NOR3_X1 i_0_2_234 (.A1(n_0_2_120), .A2(P[0]), .A3(n_0_2_104), .ZN(n_0_2_103));
   INV_X1 i_0_2_235 (.A(n_0_2_105), .ZN(n_0_2_104));
   NOR2_X1 i_0_2_236 (.A1(n_0_2_107), .A2(n_0_96), .ZN(n_0_2_105));
   OR2_X1 i_0_2_237 (.A1(reset), .A2(load), .ZN(n_0_96));
   INV_X1 i_0_2_238 (.A(n_0_2_107), .ZN(n_0_2_106));
   NOR2_X1 i_0_2_239 (.A1(n_0_2_113), .A2(n_0_2_108), .ZN(n_0_2_107));
   NAND4_X1 i_0_2_240 (.A1(n_0_2_112), .A2(n_0_2_111), .A3(n_0_2_110), .A4(
      n_0_2_109), .ZN(n_0_2_108));
   NOR4_X1 i_0_2_241 (.A1(Count[23]), .A2(Count[22]), .A3(Count[21]), .A4(
      Count[20]), .ZN(n_0_2_109));
   NOR4_X1 i_0_2_242 (.A1(Count[19]), .A2(Count[18]), .A3(Count[17]), .A4(
      Count[16]), .ZN(n_0_2_110));
   NOR4_X1 i_0_2_243 (.A1(Count[31]), .A2(Count[30]), .A3(Count[29]), .A4(
      Count[28]), .ZN(n_0_2_111));
   NOR4_X1 i_0_2_244 (.A1(Count[27]), .A2(Count[26]), .A3(Count[25]), .A4(
      Count[24]), .ZN(n_0_2_112));
   NAND4_X1 i_0_2_245 (.A1(n_0_2_117), .A2(n_0_2_116), .A3(n_0_2_115), .A4(
      n_0_2_114), .ZN(n_0_2_113));
   NOR4_X1 i_0_2_246 (.A1(Count[7]), .A2(Count[6]), .A3(Count[5]), .A4(Count[4]), 
      .ZN(n_0_2_114));
   NOR4_X1 i_0_2_247 (.A1(Count[3]), .A2(Count[2]), .A3(Count[1]), .A4(Count[0]), 
      .ZN(n_0_2_115));
   NOR4_X1 i_0_2_248 (.A1(Count[15]), .A2(Count[14]), .A3(Count[13]), .A4(
      Count[12]), .ZN(n_0_2_116));
   NOR4_X1 i_0_2_249 (.A1(Count[11]), .A2(Count[10]), .A3(Count[9]), .A4(
      Count[8]), .ZN(n_0_2_117));
   INV_X1 i_0_2_250 (.A(reset), .ZN(n_0_2_118));
   INV_X1 i_0_2_251 (.A(P[0]), .ZN(n_0_2_119));
   INV_X1 i_0_2_252 (.A(Q_minus_one), .ZN(n_0_2_120));
   DFF_X1 Q_minus_one_reg (.D(n_0_100), .CK(clk), .Q(Q_minus_one), .QN());
   MUX2_X1 Q_minus_one_reg_enable_mux_0 (.A(Q_minus_one), .B(n_0_97), .S(n_0_230), 
      .Z(n_0_100));
   CLKGATE_X1 clk_gate_Count_reg (.CK(clk), .E(n_0_165), .GCK(n_0_98));
   DFF_X1 \Count_reg[31]  (.D(n_0_229), .CK(n_0_98), .Q(Count[31]), .QN());
   DFF_X1 \Count_reg[30]  (.D(n_0_228), .CK(n_0_98), .Q(Count[30]), .QN());
   DFF_X1 \Count_reg[29]  (.D(n_0_227), .CK(n_0_98), .Q(Count[29]), .QN());
   DFF_X1 \Count_reg[28]  (.D(n_0_226), .CK(n_0_98), .Q(Count[28]), .QN());
   DFF_X1 \Count_reg[27]  (.D(n_0_225), .CK(n_0_98), .Q(Count[27]), .QN());
   DFF_X1 \Count_reg[26]  (.D(n_0_224), .CK(n_0_98), .Q(Count[26]), .QN());
   DFF_X1 \Count_reg[25]  (.D(n_0_223), .CK(n_0_98), .Q(Count[25]), .QN());
   DFF_X1 \Count_reg[24]  (.D(n_0_222), .CK(n_0_98), .Q(Count[24]), .QN());
   DFF_X1 \Count_reg[23]  (.D(n_0_221), .CK(n_0_98), .Q(Count[23]), .QN());
   DFF_X1 \Count_reg[22]  (.D(n_0_220), .CK(n_0_98), .Q(Count[22]), .QN());
   DFF_X1 \Count_reg[21]  (.D(n_0_219), .CK(n_0_98), .Q(Count[21]), .QN());
   DFF_X1 \Count_reg[20]  (.D(n_0_218), .CK(n_0_98), .Q(Count[20]), .QN());
   DFF_X1 \Count_reg[19]  (.D(n_0_217), .CK(n_0_98), .Q(Count[19]), .QN());
   DFF_X1 \Count_reg[18]  (.D(n_0_216), .CK(n_0_98), .Q(Count[18]), .QN());
   DFF_X1 \Count_reg[17]  (.D(n_0_215), .CK(n_0_98), .Q(Count[17]), .QN());
   DFF_X1 \Count_reg[16]  (.D(n_0_214), .CK(n_0_98), .Q(Count[16]), .QN());
   DFF_X1 \Count_reg[15]  (.D(n_0_213), .CK(n_0_98), .Q(Count[15]), .QN());
   DFF_X1 \Count_reg[14]  (.D(n_0_212), .CK(n_0_98), .Q(Count[14]), .QN());
   DFF_X1 \Count_reg[13]  (.D(n_0_211), .CK(n_0_98), .Q(Count[13]), .QN());
   DFF_X1 \Count_reg[12]  (.D(n_0_210), .CK(n_0_98), .Q(Count[12]), .QN());
   DFF_X1 \Count_reg[11]  (.D(n_0_209), .CK(n_0_98), .Q(Count[11]), .QN());
   DFF_X1 \Count_reg[10]  (.D(n_0_208), .CK(n_0_98), .Q(Count[10]), .QN());
   DFF_X1 \Count_reg[9]  (.D(n_0_207), .CK(n_0_98), .Q(Count[9]), .QN());
   DFF_X1 \Count_reg[8]  (.D(n_0_206), .CK(n_0_98), .Q(Count[8]), .QN());
   DFF_X1 \Count_reg[7]  (.D(n_0_205), .CK(n_0_98), .Q(Count[7]), .QN());
   DFF_X1 \Count_reg[6]  (.D(n_0_204), .CK(n_0_98), .Q(Count[6]), .QN());
   DFF_X1 \Count_reg[5]  (.D(n_0_203), .CK(n_0_98), .Q(Count[5]), .QN());
   DFF_X1 \Count_reg[4]  (.D(n_0_202), .CK(n_0_98), .Q(Count[4]), .QN());
   DFF_X1 \Count_reg[3]  (.D(n_0_201), .CK(n_0_98), .Q(Count[3]), .QN());
   DFF_X1 \Count_reg[2]  (.D(n_0_200), .CK(n_0_98), .Q(Count[2]), .QN());
   DFF_X1 \Count_reg[1]  (.D(n_0_199), .CK(n_0_98), .Q(Count[1]), .QN());
   DFF_X1 \Count_reg[0]  (.D(n_0_198), .CK(n_0_98), .Q(Count[0]), .QN());
   CLKGATE_X1 clk_gate_M_temp_reg (.CK(clk), .E(n_0_96), .GCK(n_0_99));
   DFF_X1 \M_temp_reg[31]  (.D(n_0_95), .CK(n_0_99), .Q(M_temp[31]), .QN());
   DFF_X1 \M_temp_reg[30]  (.D(n_0_94), .CK(n_0_99), .Q(M_temp[30]), .QN());
   DFF_X1 \M_temp_reg[29]  (.D(n_0_93), .CK(n_0_99), .Q(M_temp[29]), .QN());
   DFF_X1 \M_temp_reg[28]  (.D(n_0_92), .CK(n_0_99), .Q(M_temp[28]), .QN());
   DFF_X1 \M_temp_reg[27]  (.D(n_0_91), .CK(n_0_99), .Q(M_temp[27]), .QN());
   DFF_X1 \M_temp_reg[26]  (.D(n_0_90), .CK(n_0_99), .Q(M_temp[26]), .QN());
   DFF_X1 \M_temp_reg[25]  (.D(n_0_89), .CK(n_0_99), .Q(M_temp[25]), .QN());
   DFF_X1 \M_temp_reg[24]  (.D(n_0_88), .CK(n_0_99), .Q(M_temp[24]), .QN());
   DFF_X1 \M_temp_reg[23]  (.D(n_0_87), .CK(n_0_99), .Q(M_temp[23]), .QN());
   DFF_X1 \M_temp_reg[22]  (.D(n_0_86), .CK(n_0_99), .Q(M_temp[22]), .QN());
   DFF_X1 \M_temp_reg[21]  (.D(n_0_85), .CK(n_0_99), .Q(M_temp[21]), .QN());
   DFF_X1 \M_temp_reg[20]  (.D(n_0_84), .CK(n_0_99), .Q(M_temp[20]), .QN());
   DFF_X1 \M_temp_reg[19]  (.D(n_0_83), .CK(n_0_99), .Q(M_temp[19]), .QN());
   DFF_X1 \M_temp_reg[18]  (.D(n_0_82), .CK(n_0_99), .Q(M_temp[18]), .QN());
   DFF_X1 \M_temp_reg[17]  (.D(n_0_81), .CK(n_0_99), .Q(M_temp[17]), .QN());
   DFF_X1 \M_temp_reg[16]  (.D(n_0_80), .CK(n_0_99), .Q(M_temp[16]), .QN());
   DFF_X1 \M_temp_reg[15]  (.D(n_0_79), .CK(n_0_99), .Q(M_temp[15]), .QN());
   DFF_X1 \M_temp_reg[14]  (.D(n_0_78), .CK(n_0_99), .Q(M_temp[14]), .QN());
   DFF_X1 \M_temp_reg[13]  (.D(n_0_77), .CK(n_0_99), .Q(M_temp[13]), .QN());
   DFF_X1 \M_temp_reg[12]  (.D(n_0_76), .CK(n_0_99), .Q(M_temp[12]), .QN());
   DFF_X1 \M_temp_reg[11]  (.D(n_0_75), .CK(n_0_99), .Q(M_temp[11]), .QN());
   DFF_X1 \M_temp_reg[10]  (.D(n_0_74), .CK(n_0_99), .Q(M_temp[10]), .QN());
   DFF_X1 \M_temp_reg[9]  (.D(n_0_73), .CK(n_0_99), .Q(M_temp[9]), .QN());
   DFF_X1 \M_temp_reg[8]  (.D(n_0_72), .CK(n_0_99), .Q(M_temp[8]), .QN());
   DFF_X1 \M_temp_reg[7]  (.D(n_0_71), .CK(n_0_99), .Q(M_temp[7]), .QN());
   DFF_X1 \M_temp_reg[6]  (.D(n_0_70), .CK(n_0_99), .Q(M_temp[6]), .QN());
   DFF_X1 \M_temp_reg[5]  (.D(n_0_69), .CK(n_0_99), .Q(M_temp[5]), .QN());
   DFF_X1 \M_temp_reg[4]  (.D(n_0_68), .CK(n_0_99), .Q(M_temp[4]), .QN());
   DFF_X1 \M_temp_reg[3]  (.D(n_0_67), .CK(n_0_99), .Q(M_temp[3]), .QN());
   DFF_X1 \M_temp_reg[2]  (.D(n_0_66), .CK(n_0_99), .Q(M_temp[2]), .QN());
   DFF_X1 \M_temp_reg[1]  (.D(n_0_65), .CK(n_0_99), .Q(M_temp[1]), .QN());
   DFF_X1 \M_temp_reg[0]  (.D(n_0_64), .CK(n_0_99), .Q(M_temp[0]), .QN());
   DFF_X1 \P_reg[1]  (.D(n_0_102), .CK(clk), .Q(P[1]), .QN());
   DFF_X1 \P_reg[2]  (.D(n_0_103), .CK(clk), .Q(P[2]), .QN());
   DFF_X1 \P_reg[3]  (.D(n_0_104), .CK(clk), .Q(P[3]), .QN());
   DFF_X1 \P_reg[4]  (.D(n_0_105), .CK(clk), .Q(P[4]), .QN());
   DFF_X1 \P_reg[5]  (.D(n_0_106), .CK(clk), .Q(P[5]), .QN());
   DFF_X1 \P_reg[6]  (.D(n_0_107), .CK(clk), .Q(P[6]), .QN());
   DFF_X1 \P_reg[7]  (.D(n_0_108), .CK(clk), .Q(P[7]), .QN());
   DFF_X1 \P_reg[8]  (.D(n_0_109), .CK(clk), .Q(P[8]), .QN());
   DFF_X1 \P_reg[9]  (.D(n_0_110), .CK(clk), .Q(P[9]), .QN());
   DFF_X1 \P_reg[10]  (.D(n_0_111), .CK(clk), .Q(P[10]), .QN());
   DFF_X1 \P_reg[11]  (.D(n_0_112), .CK(clk), .Q(P[11]), .QN());
   DFF_X1 \P_reg[12]  (.D(n_0_113), .CK(clk), .Q(P[12]), .QN());
   DFF_X1 \P_reg[13]  (.D(n_0_114), .CK(clk), .Q(P[13]), .QN());
   DFF_X1 \P_reg[14]  (.D(n_0_115), .CK(clk), .Q(P[14]), .QN());
   DFF_X1 \P_reg[15]  (.D(n_0_116), .CK(clk), .Q(P[15]), .QN());
   DFF_X1 \P_reg[16]  (.D(n_0_117), .CK(clk), .Q(P[16]), .QN());
   DFF_X1 \P_reg[17]  (.D(n_0_118), .CK(clk), .Q(P[17]), .QN());
   DFF_X1 \P_reg[18]  (.D(n_0_119), .CK(clk), .Q(P[18]), .QN());
   DFF_X1 \P_reg[19]  (.D(n_0_120), .CK(clk), .Q(P[19]), .QN());
   DFF_X1 \P_reg[20]  (.D(n_0_121), .CK(clk), .Q(P[20]), .QN());
   DFF_X1 \P_reg[21]  (.D(n_0_122), .CK(clk), .Q(P[21]), .QN());
   DFF_X1 \P_reg[22]  (.D(n_0_123), .CK(clk), .Q(P[22]), .QN());
   DFF_X1 \P_reg[23]  (.D(n_0_124), .CK(clk), .Q(P[23]), .QN());
   DFF_X1 \P_reg[24]  (.D(n_0_125), .CK(clk), .Q(P[24]), .QN());
   DFF_X1 \P_reg[25]  (.D(n_0_126), .CK(clk), .Q(P[25]), .QN());
   DFF_X1 \P_reg[26]  (.D(n_0_127), .CK(clk), .Q(P[26]), .QN());
   DFF_X1 \P_reg[27]  (.D(n_0_128), .CK(clk), .Q(P[27]), .QN());
   DFF_X1 \P_reg[28]  (.D(n_0_129), .CK(clk), .Q(P[28]), .QN());
   DFF_X1 \P_reg[29]  (.D(n_0_130), .CK(clk), .Q(P[29]), .QN());
   DFF_X1 \P_reg[30]  (.D(n_0_131), .CK(clk), .Q(P[30]), .QN());
   DFF_X1 \P_reg[31]  (.D(n_0_132), .CK(clk), .Q(P[31]), .QN());
   DFF_X1 \P_reg[32]  (.D(n_0_133), .CK(clk), .Q(P[32]), .QN());
   DFF_X1 \P_reg[33]  (.D(n_0_134), .CK(clk), .Q(P[33]), .QN());
   DFF_X1 \P_reg[34]  (.D(n_0_135), .CK(clk), .Q(P[34]), .QN());
   DFF_X1 \P_reg[35]  (.D(n_0_136), .CK(clk), .Q(P[35]), .QN());
   DFF_X1 \P_reg[36]  (.D(n_0_137), .CK(clk), .Q(P[36]), .QN());
   DFF_X1 \P_reg[37]  (.D(n_0_138), .CK(clk), .Q(P[37]), .QN());
   DFF_X1 \P_reg[38]  (.D(n_0_139), .CK(clk), .Q(P[38]), .QN());
   DFF_X1 \P_reg[39]  (.D(n_0_140), .CK(clk), .Q(P[39]), .QN());
   DFF_X1 \P_reg[40]  (.D(n_0_141), .CK(clk), .Q(P[40]), .QN());
   DFF_X1 \P_reg[41]  (.D(n_0_142), .CK(clk), .Q(P[41]), .QN());
   DFF_X1 \P_reg[42]  (.D(n_0_143), .CK(clk), .Q(P[42]), .QN());
   DFF_X1 \P_reg[43]  (.D(n_0_144), .CK(clk), .Q(P[43]), .QN());
   DFF_X1 \P_reg[44]  (.D(n_0_145), .CK(clk), .Q(P[44]), .QN());
   DFF_X1 \P_reg[45]  (.D(n_0_146), .CK(clk), .Q(P[45]), .QN());
   DFF_X1 \P_reg[46]  (.D(n_0_147), .CK(clk), .Q(P[46]), .QN());
   DFF_X1 \P_reg[47]  (.D(n_0_148), .CK(clk), .Q(P[47]), .QN());
   DFF_X1 \P_reg[48]  (.D(n_0_149), .CK(clk), .Q(P[48]), .QN());
   DFF_X1 \P_reg[49]  (.D(n_0_150), .CK(clk), .Q(P[49]), .QN());
   DFF_X1 \P_reg[50]  (.D(n_0_151), .CK(clk), .Q(P[50]), .QN());
   DFF_X1 \P_reg[51]  (.D(n_0_152), .CK(clk), .Q(P[51]), .QN());
   DFF_X1 \P_reg[52]  (.D(n_0_153), .CK(clk), .Q(P[52]), .QN());
   DFF_X1 \P_reg[53]  (.D(n_0_154), .CK(clk), .Q(P[53]), .QN());
   DFF_X1 \P_reg[54]  (.D(n_0_155), .CK(clk), .Q(P[54]), .QN());
   DFF_X1 \P_reg[55]  (.D(n_0_156), .CK(clk), .Q(P[55]), .QN());
   DFF_X1 \P_reg[56]  (.D(n_0_157), .CK(clk), .Q(P[56]), .QN());
   DFF_X1 \P_reg[57]  (.D(n_0_158), .CK(clk), .Q(P[57]), .QN());
   DFF_X1 \P_reg[58]  (.D(n_0_159), .CK(clk), .Q(P[58]), .QN());
   DFF_X1 \P_reg[59]  (.D(n_0_160), .CK(clk), .Q(P[59]), .QN());
   DFF_X1 \P_reg[60]  (.D(n_0_161), .CK(clk), .Q(P[60]), .QN());
   DFF_X1 \P_reg[61]  (.D(n_0_162), .CK(clk), .Q(P[61]), .QN());
   DFF_X1 \P_reg[62]  (.D(n_0_163), .CK(clk), .Q(P[62]), .QN());
   DFF_X1 \P_reg[0]  (.D(n_0_101), .CK(clk), .Q(P[0]), .QN());
   DFF_X1 \P_reg[63]  (.D(n_0_164), .CK(clk), .Q(P[63]), .QN());
endmodule
