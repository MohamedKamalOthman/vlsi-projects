/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Dec 17 15:17:10 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2682476044 */

module n_case(A, B, S, outA, outB, enable);
   input [31:0]A;
   input [31:0]B;
   output [31:0]S;
   output [2:0]outA;
   output [2:0]outB;
   output enable;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_3_0;
   wire n_3_1;
   wire n_3_2;
   wire n_3_3;
   wire n_3_4;
   wire n_3_5;
   wire n_3_6;
   wire n_4_0;
   wire n_4_1;
   wire n_4_2;
   wire n_4_3;
   wire n_4_4;
   wire n_4_5;
   wire n_6_0;
   wire n_6_1;
   wire n_6_2;
   wire n_6_3;
   wire n_6_4;
   wire n_6_5;
   wire n_6_6;
   wire n_6_7;
   wire n_7_0;
   wire n_7_1;
   wire n_8_0;
   wire n_8_1;
   wire n_8_2;
   wire n_8_3;
   wire n_8_4;
   wire n_8_5;
   wire n_8_6;
   wire n_9_0;
   wire n_9_1;
   wire n_9_2;
   wire n_9_3;
   wire n_9_4;
   wire n_11_0;
   wire n_11_1;
   wire n_11_2;
   wire n_11_3;
   wire n_11_4;
   wire n_11_5;
   wire n_11_6;
   wire n_12_0;
   wire n_12_1;
   wire n_12_2;
   wire n_12_3;
   wire n_12_4;
   wire n_12_5;
   wire n_14_0;
   wire n_14_1;
   wire n_14_2;
   wire n_14_3;
   wire n_14_4;
   wire n_14_5;
   wire n_14_6;
   wire n_14_7;
   wire n_15_0;
   wire n_15_1;
   wire n_20_0;
   wire n_20_1;
   wire n_20_2;
   wire n_20_3;

   assign S[30] = S[23];
   assign S[29] = S[23];
   assign S[28] = S[23];
   assign S[27] = S[23];
   assign S[26] = S[23];
   assign S[25] = S[23];
   assign S[24] = S[23];
   assign S[22] = S[0];
   assign S[21] = S[0];
   assign S[20] = S[0];
   assign S[19] = S[0];
   assign S[18] = S[0];
   assign S[17] = S[0];
   assign S[16] = S[0];
   assign S[15] = S[0];
   assign S[14] = S[0];
   assign S[13] = S[0];
   assign S[12] = S[0];
   assign S[11] = S[0];
   assign S[10] = S[0];
   assign S[9] = S[0];
   assign S[8] = S[0];
   assign S[7] = S[0];
   assign S[6] = S[0];
   assign S[5] = S[0];
   assign S[4] = S[0];
   assign S[3] = S[0];
   assign S[2] = S[0];
   assign S[1] = S[0];

   NOR4_X1 i_0_0 (.A1(B[7]), .A2(B[8]), .A3(B[9]), .A4(B[10]), .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(B[11]), .A2(B[12]), .A3(B[13]), .A4(B[14]), .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(B[15]), .A2(B[16]), .A3(B[17]), .A4(B[18]), .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(B[19]), .A2(B[20]), .A3(B[21]), .A4(B[22]), .ZN(n_0_3));
   NAND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(n_0_4));
   NOR4_X1 i_0_5 (.A1(n_0_4), .A2(B[4]), .A3(B[5]), .A4(B[6]), .ZN(n_0_5));
   NOR4_X1 i_0_6 (.A1(B[0]), .A2(B[1]), .A3(B[2]), .A4(B[3]), .ZN(n_0_6));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_6), .ZN(n_0));
   OR4_X1 i_1_0 (.A1(B[27]), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_1_0));
   OR4_X1 i_1_1 (.A1(n_1_0), .A2(B[24]), .A3(B[25]), .A4(B[26]), .ZN(n_1_1));
   NOR2_X1 i_1_2 (.A1(n_1_1), .A2(B[23]), .ZN(n_1));
   AND4_X1 i_1_3 (.A1(B[27]), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_1_2));
   NAND4_X1 i_1_4 (.A1(n_1_2), .A2(B[24]), .A3(B[25]), .A4(B[26]), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(B[23]), .ZN(n_1_4));
   NOR2_X1 i_1_6 (.A1(n_1_3), .A2(n_1_4), .ZN(n_2));
   AND2_X1 i_2_0 (.A1(n_2), .A2(n_0), .ZN(n_3));
   NOR4_X1 i_3_0 (.A1(B[7]), .A2(B[8]), .A3(B[9]), .A4(B[10]), .ZN(n_3_0));
   NOR4_X1 i_3_1 (.A1(B[11]), .A2(B[12]), .A3(B[13]), .A4(B[14]), .ZN(n_3_1));
   NOR4_X1 i_3_2 (.A1(B[15]), .A2(B[16]), .A3(B[17]), .A4(B[18]), .ZN(n_3_2));
   NOR4_X1 i_3_3 (.A1(B[19]), .A2(B[20]), .A3(B[21]), .A4(B[22]), .ZN(n_3_3));
   NAND4_X1 i_3_4 (.A1(n_3_0), .A2(n_3_1), .A3(n_3_2), .A4(n_3_3), .ZN(n_3_4));
   NOR4_X1 i_3_5 (.A1(n_3_4), .A2(B[4]), .A3(B[5]), .A4(B[6]), .ZN(n_3_5));
   NOR4_X1 i_3_6 (.A1(B[0]), .A2(B[1]), .A3(B[2]), .A4(B[3]), .ZN(n_3_6));
   AND2_X1 i_3_7 (.A1(n_3_5), .A2(n_3_6), .ZN(n_4));
   AND2_X1 i_4_0 (.A1(n_2), .A2(n_4), .ZN(n_5));
   INV_X1 i_4_1 (.A(n_0), .ZN(n_4_0));
   AND4_X1 i_4_2 (.A1(B[27]), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_4_1));
   AND4_X1 i_4_3 (.A1(n_4_1), .A2(B[24]), .A3(B[25]), .A4(B[26]), .ZN(n_4_2));
   OR4_X1 i_4_4 (.A1(B[27]), .A2(B[28]), .A3(B[29]), .A4(B[30]), .ZN(n_4_3));
   NOR4_X1 i_4_5 (.A1(n_4_3), .A2(B[24]), .A3(B[25]), .A4(B[26]), .ZN(n_4_4));
   INV_X1 i_4_6 (.A(B[23]), .ZN(n_4_5));
   AOI221_X1 i_4_7 (.A(n_4_0), .B1(n_4_2), .B2(B[23]), .C1(n_4_4), .C2(n_4_5), 
      .ZN(n_6));
   AND2_X1 i_5_0 (.A1(n_1), .A2(n_0), .ZN(n_7));
   AND2_X1 i_5_1 (.A1(n_1), .A2(n_4), .ZN(n_8));
   NOR2_X1 i_6_0 (.A1(n_5), .A2(n_6), .ZN(n_6_0));
   INV_X1 i_6_1 (.A(n_3), .ZN(n_6_1));
   AOI21_X1 i_6_2 (.A(n_6), .B1(n_6_0), .B2(n_6_1), .ZN(n_6_2));
   OR2_X1 i_6_3 (.A1(n_7), .A2(n_8), .ZN(n_6_3));
   INV_X1 i_6_4 (.A(n_7), .ZN(n_6_4));
   OAI22_X1 i_6_5 (.A1(n_6_2), .A2(n_6_3), .B1(n_8), .B2(n_6_4), .ZN(outB[0]));
   INV_X1 i_6_6 (.A(n_6_0), .ZN(n_6_5));
   INV_X1 i_6_7 (.A(n_6), .ZN(n_6_6));
   AOI21_X1 i_6_8 (.A(n_6_3), .B1(n_6_5), .B2(n_6_6), .ZN(outB[1]));
   AOI21_X1 i_6_9 (.A(n_5), .B1(n_6_0), .B2(n_3), .ZN(n_6_7));
   NOR2_X1 i_6_10 (.A1(n_6_7), .A2(n_6_3), .ZN(outB[2]));
   INV_X1 i_7_0 (.A(outB[2]), .ZN(n_7_0));
   INV_X1 i_7_1 (.A(outB[1]), .ZN(n_7_1));
   NOR3_X1 i_7_2 (.A1(n_7_0), .A2(n_7_1), .A3(outB[0]), .ZN(n_9));
   NOR3_X1 i_7_3 (.A1(outB[0]), .A2(outB[1]), .A3(outB[2]), .ZN(n_10));
   NOR3_X1 i_7_4 (.A1(n_7_0), .A2(outB[0]), .A3(outB[1]), .ZN(n_11));
   NOR4_X1 i_8_0 (.A1(A[7]), .A2(A[8]), .A3(A[9]), .A4(A[10]), .ZN(n_8_0));
   NOR4_X1 i_8_1 (.A1(A[11]), .A2(A[12]), .A3(A[13]), .A4(A[14]), .ZN(n_8_1));
   NOR4_X1 i_8_2 (.A1(A[15]), .A2(A[16]), .A3(A[17]), .A4(A[18]), .ZN(n_8_2));
   NOR4_X1 i_8_3 (.A1(A[19]), .A2(A[20]), .A3(A[21]), .A4(A[22]), .ZN(n_8_3));
   NAND4_X1 i_8_4 (.A1(n_8_0), .A2(n_8_1), .A3(n_8_2), .A4(n_8_3), .ZN(n_8_4));
   NOR4_X1 i_8_5 (.A1(n_8_4), .A2(A[4]), .A3(A[5]), .A4(A[6]), .ZN(n_8_5));
   NOR4_X1 i_8_6 (.A1(A[0]), .A2(A[1]), .A3(A[2]), .A4(A[3]), .ZN(n_8_6));
   NAND2_X1 i_8_7 (.A1(n_8_5), .A2(n_8_6), .ZN(n_12));
   OR4_X1 i_9_0 (.A1(A[27]), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_9_0));
   OR4_X1 i_9_1 (.A1(n_9_0), .A2(A[24]), .A3(A[25]), .A4(A[26]), .ZN(n_9_1));
   NOR2_X1 i_9_2 (.A1(n_9_1), .A2(A[23]), .ZN(n_13));
   AND4_X1 i_9_3 (.A1(A[27]), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_9_2));
   NAND4_X1 i_9_4 (.A1(n_9_2), .A2(A[24]), .A3(A[25]), .A4(A[26]), .ZN(n_9_3));
   INV_X1 i_9_5 (.A(A[23]), .ZN(n_9_4));
   NOR2_X1 i_9_6 (.A1(n_9_3), .A2(n_9_4), .ZN(n_14));
   AND2_X1 i_10_0 (.A1(n_14), .A2(n_12), .ZN(n_15));
   NOR4_X1 i_11_0 (.A1(A[7]), .A2(A[8]), .A3(A[9]), .A4(A[10]), .ZN(n_11_0));
   NOR4_X1 i_11_1 (.A1(A[11]), .A2(A[12]), .A3(A[13]), .A4(A[14]), .ZN(n_11_1));
   NOR4_X1 i_11_2 (.A1(A[15]), .A2(A[16]), .A3(A[17]), .A4(A[18]), .ZN(n_11_2));
   NOR4_X1 i_11_3 (.A1(A[19]), .A2(A[20]), .A3(A[21]), .A4(A[22]), .ZN(n_11_3));
   NAND4_X1 i_11_4 (.A1(n_11_0), .A2(n_11_1), .A3(n_11_2), .A4(n_11_3), .ZN(
      n_11_4));
   NOR4_X1 i_11_5 (.A1(n_11_4), .A2(A[4]), .A3(A[5]), .A4(A[6]), .ZN(n_11_5));
   NOR4_X1 i_11_6 (.A1(A[0]), .A2(A[1]), .A3(A[2]), .A4(A[3]), .ZN(n_11_6));
   AND2_X1 i_11_7 (.A1(n_11_5), .A2(n_11_6), .ZN(n_16));
   AND2_X1 i_12_0 (.A1(n_14), .A2(n_16), .ZN(n_17));
   INV_X1 i_12_1 (.A(n_12), .ZN(n_12_0));
   AND4_X1 i_12_2 (.A1(A[27]), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_12_1));
   AND4_X1 i_12_3 (.A1(n_12_1), .A2(A[24]), .A3(A[25]), .A4(A[26]), .ZN(n_12_2));
   OR4_X1 i_12_4 (.A1(A[27]), .A2(A[28]), .A3(A[29]), .A4(A[30]), .ZN(n_12_3));
   NOR4_X1 i_12_5 (.A1(n_12_3), .A2(A[24]), .A3(A[25]), .A4(A[26]), .ZN(n_12_4));
   INV_X1 i_12_6 (.A(A[23]), .ZN(n_12_5));
   AOI221_X1 i_12_7 (.A(n_12_0), .B1(n_12_2), .B2(A[23]), .C1(n_12_4), .C2(
      n_12_5), .ZN(n_18));
   AND2_X1 i_13_0 (.A1(n_13), .A2(n_12), .ZN(n_19));
   AND2_X1 i_13_1 (.A1(n_13), .A2(n_16), .ZN(n_20));
   NOR2_X1 i_14_0 (.A1(n_17), .A2(n_18), .ZN(n_14_0));
   INV_X1 i_14_1 (.A(n_15), .ZN(n_14_1));
   AOI21_X1 i_14_2 (.A(n_18), .B1(n_14_0), .B2(n_14_1), .ZN(n_14_2));
   OR2_X1 i_14_3 (.A1(n_19), .A2(n_20), .ZN(n_14_3));
   INV_X1 i_14_4 (.A(n_19), .ZN(n_14_4));
   OAI22_X1 i_14_5 (.A1(n_14_2), .A2(n_14_3), .B1(n_20), .B2(n_14_4), .ZN(
      outA[0]));
   INV_X1 i_14_6 (.A(n_14_0), .ZN(n_14_5));
   INV_X1 i_14_7 (.A(n_18), .ZN(n_14_6));
   AOI21_X1 i_14_8 (.A(n_14_3), .B1(n_14_5), .B2(n_14_6), .ZN(outA[1]));
   AOI21_X1 i_14_9 (.A(n_17), .B1(n_14_0), .B2(n_15), .ZN(n_14_7));
   NOR2_X1 i_14_10 (.A1(n_14_7), .A2(n_14_3), .ZN(outA[2]));
   INV_X1 i_15_0 (.A(outA[2]), .ZN(n_15_0));
   INV_X1 i_15_1 (.A(outA[1]), .ZN(n_15_1));
   NOR3_X1 i_15_2 (.A1(n_15_0), .A2(n_15_1), .A3(outA[0]), .ZN(n_21));
   NOR3_X1 i_15_3 (.A1(n_15_0), .A2(outA[0]), .A3(outA[1]), .ZN(n_22));
   NOR3_X1 i_15_4 (.A1(outA[0]), .A2(outA[1]), .A3(outA[2]), .ZN(n_23));
   OR2_X1 i_16_0 (.A1(n_23), .A2(n_10), .ZN(n_24));
   OR2_X1 i_17_0 (.A1(n_22), .A2(n_11), .ZN(n_25));
   NOR2_X1 i_18_0 (.A1(n_24), .A2(n_25), .ZN(n_26));
   OR2_X1 i_18_1 (.A1(n_26), .A2(n_25), .ZN(n_27));
   XOR2_X1 i_18_2 (.A(A[31]), .B(B[31]), .Z(n_28));
   AND2_X1 i_19_0 (.A1(n_11), .A2(n_23), .ZN(n_29));
   AND2_X1 i_19_1 (.A1(n_22), .A2(n_10), .ZN(n_30));
   OR2_X1 i_19_2 (.A1(n_21), .A2(n_9), .ZN(n_31));
   NOR3_X1 i_20_0 (.A1(n_29), .A2(n_30), .A3(n_31), .ZN(n_20_0));
   NAND2_X1 i_20_1 (.A1(n_20_0), .A2(n_26), .ZN(n_20_1));
   NAND2_X1 i_20_2 (.A1(n_20_1), .A2(n_20_0), .ZN(S[0]));
   NAND2_X1 i_20_3 (.A1(n_20_0), .A2(n_27), .ZN(n_20_2));
   NAND2_X1 i_20_4 (.A1(n_20_2), .A2(n_20_0), .ZN(S[23]));
   NAND2_X1 i_20_5 (.A1(n_20_0), .A2(n_28), .ZN(n_20_3));
   NAND2_X1 i_20_6 (.A1(n_20_3), .A2(n_20_0), .ZN(S[31]));
   AND2_X1 i_21_0 (.A1(outA[0]), .A2(outB[0]), .ZN(enable));
endmodule

module zero_counter(M, Zcount);
   input [23:0]M;
   output [4:0]Zcount;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;

   AOI21_X1 i_0_0 (.A(n_0_5), .B1(n_0_0), .B2(Zcount[4]), .ZN(Zcount[0]));
   OAI21_X1 i_0_1 (.A(n_0_33), .B1(M[6]), .B2(n_0_1), .ZN(n_0_0));
   NOR2_X1 i_0_2 (.A1(M[5]), .A2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(M[4]), .A2(n_0_3), .ZN(n_0_2));
   NOR2_X1 i_0_4 (.A1(M[3]), .A2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(M[2]), .B1(n_0_32), .B2(M[0]), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(n_0_6), .B1(n_0_9), .B2(n_0_27), .ZN(n_0_5));
   AOI211_X1 i_0_7 (.A(M[15]), .B(n_0_27), .C1(n_0_7), .C2(n_0_36), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_35), .B1(M[12]), .B2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(M[11]), .B1(n_0_34), .B2(M[9]), .ZN(n_0_8));
   AOI221_X1 i_0_10 (.A(M[23]), .B1(n_0_39), .B2(M[21]), .C1(n_0_30), .C2(n_0_10), 
      .ZN(n_0_9));
   OAI21_X1 i_0_11 (.A(n_0_38), .B1(n_0_37), .B2(M[18]), .ZN(n_0_10));
   AOI21_X1 i_0_12 (.A(n_0_14), .B1(n_0_11), .B2(Zcount[4]), .ZN(Zcount[1]));
   OR3_X1 i_0_13 (.A1(M[7]), .A2(M[6]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(M[5]), .A2(M[4]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(M[3]), .A2(M[2]), .A3(n_0_23), .ZN(n_0_13));
   AOI22_X1 i_0_16 (.A1(n_0_26), .A2(n_0_17), .B1(n_0_15), .B2(n_0_27), .ZN(
      n_0_14));
   NOR3_X1 i_0_17 (.A1(M[23]), .A2(M[22]), .A3(n_0_16), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(M[21]), .A2(M[20]), .A3(n_0_29), .ZN(n_0_16));
   OAI21_X1 i_0_19 (.A(n_0_25), .B1(M[10]), .B2(M[11]), .ZN(n_0_17));
   OAI21_X1 i_0_20 (.A(n_0_18), .B1(n_0_19), .B2(Zcount[4]), .ZN(Zcount[2]));
   NAND3_X1 i_0_21 (.A1(Zcount[4]), .A2(n_0_22), .A3(n_0_21), .ZN(n_0_18));
   AOI22_X1 i_0_22 (.A1(n_0_26), .A2(n_0_25), .B1(n_0_30), .B2(n_0_27), .ZN(
      n_0_19));
   OAI22_X1 i_0_23 (.A1(n_0_22), .A2(n_0_20), .B1(n_0_27), .B2(Zcount[4]), 
      .ZN(Zcount[3]));
   NAND2_X1 i_0_24 (.A1(Zcount[4]), .A2(n_0_21), .ZN(n_0_20));
   NOR4_X1 i_0_25 (.A1(M[7]), .A2(M[6]), .A3(M[5]), .A4(M[4]), .ZN(n_0_21));
   NAND2_X1 i_0_26 (.A1(n_0_24), .A2(n_0_23), .ZN(n_0_22));
   NOR2_X1 i_0_27 (.A1(M[1]), .A2(M[0]), .ZN(n_0_23));
   NOR2_X1 i_0_28 (.A1(M[3]), .A2(M[2]), .ZN(n_0_24));
   AND3_X1 i_0_29 (.A1(n_0_31), .A2(n_0_26), .A3(n_0_25), .ZN(Zcount[4]));
   NOR2_X1 i_0_30 (.A1(M[13]), .A2(M[12]), .ZN(n_0_25));
   NOR3_X1 i_0_31 (.A1(n_0_27), .A2(M[14]), .A3(M[15]), .ZN(n_0_26));
   NAND3_X1 i_0_32 (.A1(n_0_30), .A2(n_0_29), .A3(n_0_28), .ZN(n_0_27));
   NOR2_X1 i_0_33 (.A1(M[17]), .A2(M[16]), .ZN(n_0_28));
   NOR2_X1 i_0_34 (.A1(M[19]), .A2(M[18]), .ZN(n_0_29));
   NOR4_X1 i_0_35 (.A1(M[23]), .A2(M[22]), .A3(M[21]), .A4(M[20]), .ZN(n_0_30));
   NOR4_X1 i_0_36 (.A1(M[11]), .A2(M[10]), .A3(M[9]), .A4(M[8]), .ZN(n_0_31));
   INV_X1 i_0_37 (.A(M[1]), .ZN(n_0_32));
   INV_X1 i_0_38 (.A(M[7]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(M[10]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(M[13]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(M[14]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(M[17]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(M[19]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(M[22]), .ZN(n_0_39));
endmodule

module datapath(shamt, subn, Nb);
   input [4:0]shamt;
   input [23:0]subn;
   output [23:0]Nb;

   NOR2_X1 i_0 (.A1(n_1), .A2(shamt[4]), .ZN(n_0));
   INV_X1 i_1 (.A(subn[0]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(n_3), .A2(shamt[4]), .ZN(n_2));
   INV_X1 i_3 (.A(subn[1]), .ZN(n_3));
   NOR2_X1 i_4 (.A1(n_5), .A2(shamt[4]), .ZN(n_4));
   INV_X1 i_5 (.A(subn[2]), .ZN(n_5));
   NOR2_X1 i_6 (.A1(n_7), .A2(shamt[4]), .ZN(n_6));
   INV_X1 i_7 (.A(subn[3]), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_9), .A2(shamt[4]), .ZN(n_8));
   INV_X1 i_9 (.A(subn[4]), .ZN(n_9));
   NOR2_X1 i_10 (.A1(n_11), .A2(shamt[4]), .ZN(n_10));
   INV_X1 i_11 (.A(subn[5]), .ZN(n_11));
   NOR2_X1 i_12 (.A1(n_13), .A2(shamt[4]), .ZN(n_12));
   INV_X1 i_13 (.A(subn[6]), .ZN(n_13));
   NOR2_X1 i_14 (.A1(n_15), .A2(shamt[4]), .ZN(n_14));
   INV_X1 i_15 (.A(subn[7]), .ZN(n_15));
   NOR2_X1 i_16 (.A1(n_17), .A2(shamt[4]), .ZN(n_16));
   INV_X1 i_17 (.A(subn[8]), .ZN(n_17));
   NOR2_X1 i_18 (.A1(n_19), .A2(shamt[4]), .ZN(n_18));
   INV_X1 i_19 (.A(subn[9]), .ZN(n_19));
   NOR2_X1 i_20 (.A1(n_21), .A2(shamt[4]), .ZN(n_20));
   INV_X1 i_21 (.A(subn[10]), .ZN(n_21));
   NOR2_X1 i_22 (.A1(n_23), .A2(shamt[4]), .ZN(n_22));
   INV_X1 i_23 (.A(subn[11]), .ZN(n_23));
   NOR2_X1 i_24 (.A1(n_25), .A2(shamt[4]), .ZN(n_24));
   INV_X1 i_25 (.A(subn[12]), .ZN(n_25));
   NOR2_X1 i_26 (.A1(n_27), .A2(shamt[4]), .ZN(n_26));
   INV_X1 i_27 (.A(subn[13]), .ZN(n_27));
   NOR2_X1 i_28 (.A1(n_29), .A2(shamt[4]), .ZN(n_28));
   INV_X1 i_29 (.A(subn[14]), .ZN(n_29));
   NOR2_X1 i_30 (.A1(n_31), .A2(shamt[4]), .ZN(n_30));
   INV_X1 i_31 (.A(subn[15]), .ZN(n_31));
   MUX2_X1 i_32 (.A(subn[16]), .B(subn[0]), .S(shamt[4]), .Z(n_32));
   MUX2_X1 i_33 (.A(subn[17]), .B(subn[1]), .S(shamt[4]), .Z(n_33));
   MUX2_X1 i_34 (.A(subn[18]), .B(subn[2]), .S(shamt[4]), .Z(n_34));
   MUX2_X1 i_35 (.A(subn[19]), .B(subn[3]), .S(shamt[4]), .Z(n_35));
   MUX2_X1 i_36 (.A(subn[20]), .B(subn[4]), .S(shamt[4]), .Z(n_36));
   MUX2_X1 i_37 (.A(subn[21]), .B(subn[5]), .S(shamt[4]), .Z(n_37));
   MUX2_X1 i_38 (.A(subn[22]), .B(subn[6]), .S(shamt[4]), .Z(n_38));
   MUX2_X1 i_39 (.A(subn[23]), .B(subn[7]), .S(shamt[4]), .Z(n_39));
   NOR2_X1 i_40 (.A1(n_41), .A2(shamt[3]), .ZN(n_40));
   INV_X1 i_41 (.A(n_0), .ZN(n_41));
   NOR2_X1 i_42 (.A1(n_43), .A2(shamt[3]), .ZN(n_42));
   INV_X1 i_43 (.A(n_2), .ZN(n_43));
   NOR2_X1 i_44 (.A1(n_45), .A2(shamt[3]), .ZN(n_44));
   INV_X1 i_45 (.A(n_4), .ZN(n_45));
   NOR2_X1 i_46 (.A1(n_47), .A2(shamt[3]), .ZN(n_46));
   INV_X1 i_47 (.A(n_6), .ZN(n_47));
   NOR2_X1 i_48 (.A1(n_49), .A2(shamt[3]), .ZN(n_48));
   INV_X1 i_49 (.A(n_8), .ZN(n_49));
   NOR2_X1 i_50 (.A1(n_51), .A2(shamt[3]), .ZN(n_50));
   INV_X1 i_51 (.A(n_10), .ZN(n_51));
   NOR2_X1 i_52 (.A1(n_53), .A2(shamt[3]), .ZN(n_52));
   INV_X1 i_53 (.A(n_12), .ZN(n_53));
   NOR2_X1 i_54 (.A1(n_55), .A2(shamt[3]), .ZN(n_54));
   INV_X1 i_55 (.A(n_14), .ZN(n_55));
   MUX2_X1 i_56 (.A(n_16), .B(n_0), .S(shamt[3]), .Z(n_56));
   MUX2_X1 i_57 (.A(n_18), .B(n_2), .S(shamt[3]), .Z(n_57));
   MUX2_X1 i_58 (.A(n_20), .B(n_4), .S(shamt[3]), .Z(n_58));
   MUX2_X1 i_59 (.A(n_22), .B(n_6), .S(shamt[3]), .Z(n_59));
   MUX2_X1 i_60 (.A(n_24), .B(n_8), .S(shamt[3]), .Z(n_60));
   MUX2_X1 i_61 (.A(n_26), .B(n_10), .S(shamt[3]), .Z(n_61));
   MUX2_X1 i_62 (.A(n_28), .B(n_12), .S(shamt[3]), .Z(n_62));
   MUX2_X1 i_63 (.A(n_30), .B(n_14), .S(shamt[3]), .Z(n_63));
   MUX2_X1 i_64 (.A(n_32), .B(n_16), .S(shamt[3]), .Z(n_64));
   MUX2_X1 i_65 (.A(n_33), .B(n_18), .S(shamt[3]), .Z(n_65));
   MUX2_X1 i_66 (.A(n_34), .B(n_20), .S(shamt[3]), .Z(n_66));
   MUX2_X1 i_67 (.A(n_35), .B(n_22), .S(shamt[3]), .Z(n_67));
   MUX2_X1 i_68 (.A(n_36), .B(n_24), .S(shamt[3]), .Z(n_68));
   MUX2_X1 i_69 (.A(n_37), .B(n_26), .S(shamt[3]), .Z(n_69));
   MUX2_X1 i_70 (.A(n_38), .B(n_28), .S(shamt[3]), .Z(n_70));
   MUX2_X1 i_71 (.A(n_39), .B(n_30), .S(shamt[3]), .Z(n_71));
   NOR2_X1 i_72 (.A1(n_73), .A2(shamt[2]), .ZN(n_72));
   INV_X1 i_73 (.A(n_40), .ZN(n_73));
   NOR2_X1 i_74 (.A1(n_75), .A2(shamt[2]), .ZN(n_74));
   INV_X1 i_75 (.A(n_42), .ZN(n_75));
   NOR2_X1 i_76 (.A1(n_77), .A2(shamt[2]), .ZN(n_76));
   INV_X1 i_77 (.A(n_44), .ZN(n_77));
   NOR2_X1 i_78 (.A1(n_79), .A2(shamt[2]), .ZN(n_78));
   INV_X1 i_79 (.A(n_46), .ZN(n_79));
   MUX2_X1 i_80 (.A(n_48), .B(n_40), .S(shamt[2]), .Z(n_80));
   MUX2_X1 i_81 (.A(n_50), .B(n_42), .S(shamt[2]), .Z(n_81));
   MUX2_X1 i_82 (.A(n_52), .B(n_44), .S(shamt[2]), .Z(n_82));
   MUX2_X1 i_83 (.A(n_54), .B(n_46), .S(shamt[2]), .Z(n_83));
   MUX2_X1 i_84 (.A(n_56), .B(n_48), .S(shamt[2]), .Z(n_84));
   MUX2_X1 i_85 (.A(n_57), .B(n_50), .S(shamt[2]), .Z(n_85));
   MUX2_X1 i_86 (.A(n_58), .B(n_52), .S(shamt[2]), .Z(n_86));
   MUX2_X1 i_87 (.A(n_59), .B(n_54), .S(shamt[2]), .Z(n_87));
   MUX2_X1 i_88 (.A(n_60), .B(n_56), .S(shamt[2]), .Z(n_88));
   MUX2_X1 i_89 (.A(n_61), .B(n_57), .S(shamt[2]), .Z(n_89));
   MUX2_X1 i_90 (.A(n_62), .B(n_58), .S(shamt[2]), .Z(n_90));
   MUX2_X1 i_91 (.A(n_63), .B(n_59), .S(shamt[2]), .Z(n_91));
   MUX2_X1 i_92 (.A(n_64), .B(n_60), .S(shamt[2]), .Z(n_92));
   MUX2_X1 i_93 (.A(n_65), .B(n_61), .S(shamt[2]), .Z(n_93));
   MUX2_X1 i_94 (.A(n_66), .B(n_62), .S(shamt[2]), .Z(n_94));
   MUX2_X1 i_95 (.A(n_67), .B(n_63), .S(shamt[2]), .Z(n_95));
   MUX2_X1 i_96 (.A(n_68), .B(n_64), .S(shamt[2]), .Z(n_96));
   MUX2_X1 i_97 (.A(n_69), .B(n_65), .S(shamt[2]), .Z(n_97));
   MUX2_X1 i_98 (.A(n_70), .B(n_66), .S(shamt[2]), .Z(n_98));
   MUX2_X1 i_99 (.A(n_71), .B(n_67), .S(shamt[2]), .Z(n_99));
   NOR2_X1 i_100 (.A1(n_101), .A2(shamt[1]), .ZN(n_100));
   INV_X1 i_101 (.A(n_72), .ZN(n_101));
   NOR2_X1 i_102 (.A1(n_103), .A2(shamt[1]), .ZN(n_102));
   INV_X1 i_103 (.A(n_74), .ZN(n_103));
   MUX2_X1 i_104 (.A(n_76), .B(n_72), .S(shamt[1]), .Z(n_104));
   MUX2_X1 i_105 (.A(n_78), .B(n_74), .S(shamt[1]), .Z(n_105));
   MUX2_X1 i_106 (.A(n_80), .B(n_76), .S(shamt[1]), .Z(n_106));
   MUX2_X1 i_107 (.A(n_81), .B(n_78), .S(shamt[1]), .Z(n_107));
   MUX2_X1 i_108 (.A(n_82), .B(n_80), .S(shamt[1]), .Z(n_108));
   MUX2_X1 i_109 (.A(n_83), .B(n_81), .S(shamt[1]), .Z(n_109));
   MUX2_X1 i_110 (.A(n_84), .B(n_82), .S(shamt[1]), .Z(n_110));
   MUX2_X1 i_111 (.A(n_85), .B(n_83), .S(shamt[1]), .Z(n_111));
   MUX2_X1 i_112 (.A(n_86), .B(n_84), .S(shamt[1]), .Z(n_112));
   MUX2_X1 i_113 (.A(n_87), .B(n_85), .S(shamt[1]), .Z(n_113));
   MUX2_X1 i_114 (.A(n_88), .B(n_86), .S(shamt[1]), .Z(n_114));
   MUX2_X1 i_115 (.A(n_89), .B(n_87), .S(shamt[1]), .Z(n_115));
   MUX2_X1 i_116 (.A(n_90), .B(n_88), .S(shamt[1]), .Z(n_116));
   MUX2_X1 i_117 (.A(n_91), .B(n_89), .S(shamt[1]), .Z(n_117));
   MUX2_X1 i_118 (.A(n_92), .B(n_90), .S(shamt[1]), .Z(n_118));
   MUX2_X1 i_119 (.A(n_93), .B(n_91), .S(shamt[1]), .Z(n_119));
   MUX2_X1 i_120 (.A(n_94), .B(n_92), .S(shamt[1]), .Z(n_120));
   MUX2_X1 i_121 (.A(n_95), .B(n_93), .S(shamt[1]), .Z(n_121));
   MUX2_X1 i_122 (.A(n_96), .B(n_94), .S(shamt[1]), .Z(n_122));
   MUX2_X1 i_123 (.A(n_97), .B(n_95), .S(shamt[1]), .Z(n_123));
   MUX2_X1 i_124 (.A(n_98), .B(n_96), .S(shamt[1]), .Z(n_124));
   MUX2_X1 i_125 (.A(n_99), .B(n_97), .S(shamt[1]), .Z(n_125));
   NOR2_X1 i_126 (.A1(n_126), .A2(shamt[0]), .ZN(Nb[0]));
   INV_X1 i_127 (.A(n_100), .ZN(n_126));
   MUX2_X1 i_128 (.A(n_102), .B(n_100), .S(shamt[0]), .Z(Nb[1]));
   MUX2_X1 i_129 (.A(n_104), .B(n_102), .S(shamt[0]), .Z(Nb[2]));
   MUX2_X1 i_130 (.A(n_105), .B(n_104), .S(shamt[0]), .Z(Nb[3]));
   MUX2_X1 i_131 (.A(n_106), .B(n_105), .S(shamt[0]), .Z(Nb[4]));
   MUX2_X1 i_132 (.A(n_107), .B(n_106), .S(shamt[0]), .Z(Nb[5]));
   MUX2_X1 i_133 (.A(n_108), .B(n_107), .S(shamt[0]), .Z(Nb[6]));
   MUX2_X1 i_134 (.A(n_109), .B(n_108), .S(shamt[0]), .Z(Nb[7]));
   MUX2_X1 i_135 (.A(n_110), .B(n_109), .S(shamt[0]), .Z(Nb[8]));
   MUX2_X1 i_136 (.A(n_111), .B(n_110), .S(shamt[0]), .Z(Nb[9]));
   MUX2_X1 i_137 (.A(n_112), .B(n_111), .S(shamt[0]), .Z(Nb[10]));
   MUX2_X1 i_138 (.A(n_113), .B(n_112), .S(shamt[0]), .Z(Nb[11]));
   MUX2_X1 i_139 (.A(n_114), .B(n_113), .S(shamt[0]), .Z(Nb[12]));
   MUX2_X1 i_140 (.A(n_115), .B(n_114), .S(shamt[0]), .Z(Nb[13]));
   MUX2_X1 i_141 (.A(n_116), .B(n_115), .S(shamt[0]), .Z(Nb[14]));
   MUX2_X1 i_142 (.A(n_117), .B(n_116), .S(shamt[0]), .Z(Nb[15]));
   MUX2_X1 i_143 (.A(n_118), .B(n_117), .S(shamt[0]), .Z(Nb[16]));
   MUX2_X1 i_144 (.A(n_119), .B(n_118), .S(shamt[0]), .Z(Nb[17]));
   MUX2_X1 i_145 (.A(n_120), .B(n_119), .S(shamt[0]), .Z(Nb[18]));
   MUX2_X1 i_146 (.A(n_121), .B(n_120), .S(shamt[0]), .Z(Nb[19]));
   MUX2_X1 i_147 (.A(n_122), .B(n_121), .S(shamt[0]), .Z(Nb[20]));
   MUX2_X1 i_148 (.A(n_123), .B(n_122), .S(shamt[0]), .Z(Nb[21]));
   MUX2_X1 i_149 (.A(n_124), .B(n_123), .S(shamt[0]), .Z(Nb[22]));
   MUX2_X1 i_150 (.A(n_125), .B(n_124), .S(shamt[0]), .Z(Nb[23]));
endmodule

module datapath__0_29(Nb, Na, mult_res);
   input [23:0]Nb;
   input [23:0]Na;
   output [47:0]mult_res;

   NAND2_X1 i_0 (.A1(Nb[0]), .A2(Na[1]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(Nb[0]), .A2(Na[2]), .ZN(n_1));
   NAND2_X1 i_2 (.A1(Nb[0]), .A2(Na[3]), .ZN(n_2));
   NAND2_X1 i_3 (.A1(Nb[0]), .A2(Na[4]), .ZN(n_3));
   NAND2_X1 i_4 (.A1(Nb[0]), .A2(Na[5]), .ZN(n_4));
   NAND2_X1 i_5 (.A1(Nb[0]), .A2(Na[6]), .ZN(n_5));
   NAND2_X1 i_6 (.A1(Nb[0]), .A2(Na[7]), .ZN(n_6));
   NAND2_X1 i_7 (.A1(Nb[0]), .A2(Na[8]), .ZN(n_7));
   NAND2_X1 i_8 (.A1(Nb[0]), .A2(Na[9]), .ZN(n_8));
   NAND2_X1 i_9 (.A1(Nb[0]), .A2(Na[10]), .ZN(n_9));
   NAND2_X1 i_10 (.A1(Nb[0]), .A2(Na[11]), .ZN(n_10));
   NAND2_X1 i_11 (.A1(Nb[0]), .A2(Na[12]), .ZN(n_11));
   NAND2_X1 i_12 (.A1(Nb[0]), .A2(Na[13]), .ZN(n_12));
   NAND2_X1 i_13 (.A1(Nb[0]), .A2(Na[14]), .ZN(n_13));
   NAND2_X1 i_14 (.A1(Nb[0]), .A2(Na[15]), .ZN(n_14));
   NAND2_X1 i_15 (.A1(Nb[0]), .A2(Na[16]), .ZN(n_15));
   NAND2_X1 i_16 (.A1(Nb[0]), .A2(Na[17]), .ZN(n_16));
   NAND2_X1 i_17 (.A1(Nb[0]), .A2(Na[18]), .ZN(n_17));
   NAND2_X1 i_18 (.A1(Nb[0]), .A2(Na[19]), .ZN(n_18));
   NAND2_X1 i_19 (.A1(Nb[0]), .A2(Na[20]), .ZN(n_19));
   NAND2_X1 i_20 (.A1(Nb[0]), .A2(Na[21]), .ZN(n_20));
   NAND2_X1 i_21 (.A1(Nb[0]), .A2(Na[22]), .ZN(n_21));
   NAND2_X1 i_22 (.A1(Nb[0]), .A2(Na[23]), .ZN(n_22));
   NAND2_X1 i_23 (.A1(Nb[1]), .A2(Na[0]), .ZN(n_23));
   NAND2_X1 i_24 (.A1(Nb[1]), .A2(Na[1]), .ZN(n_24));
   NAND2_X1 i_25 (.A1(Nb[1]), .A2(Na[2]), .ZN(n_25));
   NAND2_X1 i_26 (.A1(Nb[1]), .A2(Na[3]), .ZN(n_26));
   NAND2_X1 i_27 (.A1(Nb[1]), .A2(Na[4]), .ZN(n_27));
   NAND2_X1 i_28 (.A1(Nb[1]), .A2(Na[5]), .ZN(n_28));
   NAND2_X1 i_29 (.A1(Nb[1]), .A2(Na[6]), .ZN(n_29));
   NAND2_X1 i_30 (.A1(Nb[1]), .A2(Na[7]), .ZN(n_30));
   NAND2_X1 i_31 (.A1(Nb[1]), .A2(Na[8]), .ZN(n_31));
   NAND2_X1 i_32 (.A1(Nb[1]), .A2(Na[9]), .ZN(n_32));
   NAND2_X1 i_33 (.A1(Nb[1]), .A2(Na[10]), .ZN(n_33));
   NAND2_X1 i_34 (.A1(Nb[1]), .A2(Na[11]), .ZN(n_34));
   NAND2_X1 i_35 (.A1(Nb[1]), .A2(Na[12]), .ZN(n_35));
   NAND2_X1 i_36 (.A1(Nb[1]), .A2(Na[13]), .ZN(n_36));
   NAND2_X1 i_37 (.A1(Nb[1]), .A2(Na[14]), .ZN(n_37));
   NAND2_X1 i_38 (.A1(Nb[1]), .A2(Na[15]), .ZN(n_38));
   NAND2_X1 i_39 (.A1(Nb[1]), .A2(Na[16]), .ZN(n_39));
   NAND2_X1 i_40 (.A1(Nb[1]), .A2(Na[17]), .ZN(n_40));
   NAND2_X1 i_41 (.A1(Nb[1]), .A2(Na[18]), .ZN(n_41));
   NAND2_X1 i_42 (.A1(Nb[1]), .A2(Na[19]), .ZN(n_42));
   NAND2_X1 i_43 (.A1(Nb[1]), .A2(Na[20]), .ZN(n_43));
   NAND2_X1 i_44 (.A1(Nb[1]), .A2(Na[21]), .ZN(n_44));
   NAND2_X1 i_45 (.A1(Nb[1]), .A2(Na[22]), .ZN(n_45));
   NAND2_X1 i_46 (.A1(Nb[1]), .A2(Na[23]), .ZN(n_46));
   NAND2_X1 i_47 (.A1(Nb[2]), .A2(Na[0]), .ZN(n_47));
   NAND2_X1 i_48 (.A1(Nb[2]), .A2(Na[1]), .ZN(n_48));
   NAND2_X1 i_49 (.A1(Nb[2]), .A2(Na[2]), .ZN(n_49));
   NAND2_X1 i_50 (.A1(Nb[2]), .A2(Na[3]), .ZN(n_50));
   NAND2_X1 i_51 (.A1(Nb[2]), .A2(Na[4]), .ZN(n_51));
   NAND2_X1 i_52 (.A1(Nb[2]), .A2(Na[5]), .ZN(n_52));
   NAND2_X1 i_53 (.A1(Nb[2]), .A2(Na[6]), .ZN(n_53));
   NAND2_X1 i_54 (.A1(Nb[2]), .A2(Na[7]), .ZN(n_54));
   NAND2_X1 i_55 (.A1(Nb[2]), .A2(Na[8]), .ZN(n_55));
   NAND2_X1 i_56 (.A1(Nb[2]), .A2(Na[9]), .ZN(n_56));
   NAND2_X1 i_57 (.A1(Nb[2]), .A2(Na[10]), .ZN(n_57));
   NAND2_X1 i_58 (.A1(Nb[2]), .A2(Na[11]), .ZN(n_58));
   NAND2_X1 i_59 (.A1(Nb[2]), .A2(Na[12]), .ZN(n_59));
   NAND2_X1 i_60 (.A1(Nb[2]), .A2(Na[13]), .ZN(n_60));
   NAND2_X1 i_61 (.A1(Nb[2]), .A2(Na[14]), .ZN(n_61));
   NAND2_X1 i_62 (.A1(Nb[2]), .A2(Na[15]), .ZN(n_62));
   NAND2_X1 i_63 (.A1(Nb[2]), .A2(Na[16]), .ZN(n_63));
   NAND2_X1 i_64 (.A1(Nb[2]), .A2(Na[17]), .ZN(n_64));
   NAND2_X1 i_65 (.A1(Nb[2]), .A2(Na[18]), .ZN(n_65));
   NAND2_X1 i_66 (.A1(Nb[2]), .A2(Na[19]), .ZN(n_66));
   NAND2_X1 i_67 (.A1(Nb[2]), .A2(Na[20]), .ZN(n_67));
   NAND2_X1 i_68 (.A1(Nb[2]), .A2(Na[21]), .ZN(n_68));
   NAND2_X1 i_69 (.A1(Nb[2]), .A2(Na[22]), .ZN(n_69));
   NAND2_X1 i_70 (.A1(Nb[2]), .A2(Na[23]), .ZN(n_70));
   NAND2_X1 i_71 (.A1(Nb[3]), .A2(Na[0]), .ZN(n_71));
   NAND2_X1 i_72 (.A1(Nb[3]), .A2(Na[1]), .ZN(n_72));
   NAND2_X1 i_73 (.A1(Nb[3]), .A2(Na[2]), .ZN(n_73));
   NAND2_X1 i_74 (.A1(Nb[3]), .A2(Na[3]), .ZN(n_74));
   NAND2_X1 i_75 (.A1(Nb[3]), .A2(Na[4]), .ZN(n_75));
   NAND2_X1 i_76 (.A1(Nb[3]), .A2(Na[5]), .ZN(n_76));
   NAND2_X1 i_77 (.A1(Nb[3]), .A2(Na[6]), .ZN(n_77));
   NAND2_X1 i_78 (.A1(Nb[3]), .A2(Na[7]), .ZN(n_78));
   NAND2_X1 i_79 (.A1(Nb[3]), .A2(Na[8]), .ZN(n_79));
   NAND2_X1 i_80 (.A1(Nb[3]), .A2(Na[9]), .ZN(n_80));
   NAND2_X1 i_81 (.A1(Nb[3]), .A2(Na[10]), .ZN(n_81));
   NAND2_X1 i_82 (.A1(Nb[3]), .A2(Na[11]), .ZN(n_82));
   NAND2_X1 i_83 (.A1(Nb[3]), .A2(Na[12]), .ZN(n_83));
   NAND2_X1 i_84 (.A1(Nb[3]), .A2(Na[13]), .ZN(n_84));
   NAND2_X1 i_85 (.A1(Nb[3]), .A2(Na[14]), .ZN(n_85));
   NAND2_X1 i_86 (.A1(Nb[3]), .A2(Na[15]), .ZN(n_86));
   NAND2_X1 i_87 (.A1(Nb[3]), .A2(Na[16]), .ZN(n_87));
   NAND2_X1 i_88 (.A1(Nb[3]), .A2(Na[17]), .ZN(n_88));
   NAND2_X1 i_89 (.A1(Nb[3]), .A2(Na[18]), .ZN(n_89));
   NAND2_X1 i_90 (.A1(Nb[3]), .A2(Na[19]), .ZN(n_90));
   NAND2_X1 i_91 (.A1(Nb[3]), .A2(Na[20]), .ZN(n_91));
   NAND2_X1 i_92 (.A1(Nb[3]), .A2(Na[21]), .ZN(n_92));
   NAND2_X1 i_93 (.A1(Nb[3]), .A2(Na[22]), .ZN(n_93));
   NAND2_X1 i_94 (.A1(Nb[3]), .A2(Na[23]), .ZN(n_94));
   NAND2_X1 i_95 (.A1(Nb[4]), .A2(Na[0]), .ZN(n_95));
   NAND2_X1 i_96 (.A1(Nb[4]), .A2(Na[1]), .ZN(n_96));
   NAND2_X1 i_97 (.A1(Nb[4]), .A2(Na[2]), .ZN(n_97));
   NAND2_X1 i_98 (.A1(Nb[4]), .A2(Na[3]), .ZN(n_98));
   NAND2_X1 i_99 (.A1(Nb[4]), .A2(Na[4]), .ZN(n_99));
   NAND2_X1 i_100 (.A1(Nb[4]), .A2(Na[5]), .ZN(n_100));
   NAND2_X1 i_101 (.A1(Nb[4]), .A2(Na[6]), .ZN(n_101));
   NAND2_X1 i_102 (.A1(Nb[4]), .A2(Na[7]), .ZN(n_102));
   NAND2_X1 i_103 (.A1(Nb[4]), .A2(Na[8]), .ZN(n_103));
   NAND2_X1 i_104 (.A1(Nb[4]), .A2(Na[9]), .ZN(n_104));
   NAND2_X1 i_105 (.A1(Nb[4]), .A2(Na[10]), .ZN(n_105));
   NAND2_X1 i_106 (.A1(Nb[4]), .A2(Na[11]), .ZN(n_106));
   NAND2_X1 i_107 (.A1(Nb[4]), .A2(Na[12]), .ZN(n_107));
   NAND2_X1 i_108 (.A1(Nb[4]), .A2(Na[13]), .ZN(n_108));
   NAND2_X1 i_109 (.A1(Nb[4]), .A2(Na[14]), .ZN(n_109));
   NAND2_X1 i_110 (.A1(Nb[4]), .A2(Na[15]), .ZN(n_110));
   NAND2_X1 i_111 (.A1(Nb[4]), .A2(Na[16]), .ZN(n_111));
   NAND2_X1 i_112 (.A1(Nb[4]), .A2(Na[17]), .ZN(n_112));
   NAND2_X1 i_113 (.A1(Nb[4]), .A2(Na[18]), .ZN(n_113));
   NAND2_X1 i_114 (.A1(Nb[4]), .A2(Na[19]), .ZN(n_114));
   NAND2_X1 i_115 (.A1(Nb[4]), .A2(Na[20]), .ZN(n_115));
   NAND2_X1 i_116 (.A1(Nb[4]), .A2(Na[21]), .ZN(n_116));
   NAND2_X1 i_117 (.A1(Nb[4]), .A2(Na[22]), .ZN(n_117));
   NAND2_X1 i_118 (.A1(Nb[4]), .A2(Na[23]), .ZN(n_118));
   NAND2_X1 i_119 (.A1(Nb[5]), .A2(Na[0]), .ZN(n_119));
   NAND2_X1 i_120 (.A1(Nb[5]), .A2(Na[1]), .ZN(n_120));
   NAND2_X1 i_121 (.A1(Nb[5]), .A2(Na[2]), .ZN(n_121));
   NAND2_X1 i_122 (.A1(Nb[5]), .A2(Na[3]), .ZN(n_122));
   NAND2_X1 i_123 (.A1(Nb[5]), .A2(Na[4]), .ZN(n_123));
   NAND2_X1 i_124 (.A1(Nb[5]), .A2(Na[5]), .ZN(n_124));
   NAND2_X1 i_125 (.A1(Nb[5]), .A2(Na[6]), .ZN(n_125));
   NAND2_X1 i_126 (.A1(Nb[5]), .A2(Na[7]), .ZN(n_126));
   NAND2_X1 i_127 (.A1(Nb[5]), .A2(Na[8]), .ZN(n_127));
   NAND2_X1 i_128 (.A1(Nb[5]), .A2(Na[9]), .ZN(n_128));
   NAND2_X1 i_129 (.A1(Nb[5]), .A2(Na[10]), .ZN(n_129));
   NAND2_X1 i_130 (.A1(Nb[5]), .A2(Na[11]), .ZN(n_130));
   NAND2_X1 i_131 (.A1(Nb[5]), .A2(Na[12]), .ZN(n_131));
   NAND2_X1 i_132 (.A1(Nb[5]), .A2(Na[13]), .ZN(n_132));
   NAND2_X1 i_133 (.A1(Nb[5]), .A2(Na[14]), .ZN(n_133));
   NAND2_X1 i_134 (.A1(Nb[5]), .A2(Na[15]), .ZN(n_134));
   NAND2_X1 i_135 (.A1(Nb[5]), .A2(Na[16]), .ZN(n_135));
   NAND2_X1 i_136 (.A1(Nb[5]), .A2(Na[17]), .ZN(n_136));
   NAND2_X1 i_137 (.A1(Nb[5]), .A2(Na[18]), .ZN(n_137));
   NAND2_X1 i_138 (.A1(Nb[5]), .A2(Na[19]), .ZN(n_138));
   NAND2_X1 i_139 (.A1(Nb[5]), .A2(Na[20]), .ZN(n_139));
   NAND2_X1 i_140 (.A1(Nb[5]), .A2(Na[21]), .ZN(n_140));
   NAND2_X1 i_141 (.A1(Nb[5]), .A2(Na[22]), .ZN(n_141));
   NAND2_X1 i_142 (.A1(Nb[5]), .A2(Na[23]), .ZN(n_142));
   NAND2_X1 i_143 (.A1(Nb[6]), .A2(Na[0]), .ZN(n_143));
   NAND2_X1 i_144 (.A1(Nb[6]), .A2(Na[1]), .ZN(n_144));
   NAND2_X1 i_145 (.A1(Nb[6]), .A2(Na[2]), .ZN(n_145));
   NAND2_X1 i_146 (.A1(Nb[6]), .A2(Na[3]), .ZN(n_146));
   NAND2_X1 i_147 (.A1(Nb[6]), .A2(Na[4]), .ZN(n_147));
   NAND2_X1 i_148 (.A1(Nb[6]), .A2(Na[5]), .ZN(n_148));
   NAND2_X1 i_149 (.A1(Nb[6]), .A2(Na[6]), .ZN(n_149));
   NAND2_X1 i_150 (.A1(Nb[6]), .A2(Na[7]), .ZN(n_150));
   NAND2_X1 i_151 (.A1(Nb[6]), .A2(Na[8]), .ZN(n_151));
   NAND2_X1 i_152 (.A1(Nb[6]), .A2(Na[9]), .ZN(n_152));
   NAND2_X1 i_153 (.A1(Nb[6]), .A2(Na[10]), .ZN(n_153));
   NAND2_X1 i_154 (.A1(Nb[6]), .A2(Na[11]), .ZN(n_154));
   NAND2_X1 i_155 (.A1(Nb[6]), .A2(Na[12]), .ZN(n_155));
   NAND2_X1 i_156 (.A1(Nb[6]), .A2(Na[13]), .ZN(n_156));
   NAND2_X1 i_157 (.A1(Nb[6]), .A2(Na[14]), .ZN(n_157));
   NAND2_X1 i_158 (.A1(Nb[6]), .A2(Na[15]), .ZN(n_158));
   NAND2_X1 i_159 (.A1(Nb[6]), .A2(Na[16]), .ZN(n_159));
   NAND2_X1 i_160 (.A1(Nb[6]), .A2(Na[17]), .ZN(n_160));
   NAND2_X1 i_161 (.A1(Nb[6]), .A2(Na[18]), .ZN(n_161));
   NAND2_X1 i_162 (.A1(Nb[6]), .A2(Na[19]), .ZN(n_162));
   NAND2_X1 i_163 (.A1(Nb[6]), .A2(Na[20]), .ZN(n_163));
   NAND2_X1 i_164 (.A1(Nb[6]), .A2(Na[21]), .ZN(n_164));
   NAND2_X1 i_165 (.A1(Nb[6]), .A2(Na[22]), .ZN(n_165));
   NAND2_X1 i_166 (.A1(Nb[6]), .A2(Na[23]), .ZN(n_166));
   NAND2_X1 i_167 (.A1(Nb[7]), .A2(Na[0]), .ZN(n_167));
   NAND2_X1 i_168 (.A1(Nb[7]), .A2(Na[1]), .ZN(n_168));
   NAND2_X1 i_169 (.A1(Nb[7]), .A2(Na[2]), .ZN(n_169));
   NAND2_X1 i_170 (.A1(Nb[7]), .A2(Na[3]), .ZN(n_170));
   NAND2_X1 i_171 (.A1(Nb[7]), .A2(Na[4]), .ZN(n_171));
   NAND2_X1 i_172 (.A1(Nb[7]), .A2(Na[5]), .ZN(n_172));
   NAND2_X1 i_173 (.A1(Nb[7]), .A2(Na[6]), .ZN(n_173));
   NAND2_X1 i_174 (.A1(Nb[7]), .A2(Na[7]), .ZN(n_174));
   NAND2_X1 i_175 (.A1(Nb[7]), .A2(Na[8]), .ZN(n_175));
   NAND2_X1 i_176 (.A1(Nb[7]), .A2(Na[9]), .ZN(n_176));
   NAND2_X1 i_177 (.A1(Nb[7]), .A2(Na[10]), .ZN(n_177));
   NAND2_X1 i_178 (.A1(Nb[7]), .A2(Na[11]), .ZN(n_178));
   NAND2_X1 i_179 (.A1(Nb[7]), .A2(Na[12]), .ZN(n_179));
   NAND2_X1 i_180 (.A1(Nb[7]), .A2(Na[13]), .ZN(n_180));
   NAND2_X1 i_181 (.A1(Nb[7]), .A2(Na[14]), .ZN(n_181));
   NAND2_X1 i_182 (.A1(Nb[7]), .A2(Na[15]), .ZN(n_182));
   NAND2_X1 i_183 (.A1(Nb[7]), .A2(Na[16]), .ZN(n_183));
   NAND2_X1 i_184 (.A1(Nb[7]), .A2(Na[17]), .ZN(n_184));
   NAND2_X1 i_185 (.A1(Nb[7]), .A2(Na[18]), .ZN(n_185));
   NAND2_X1 i_186 (.A1(Nb[7]), .A2(Na[19]), .ZN(n_186));
   NAND2_X1 i_187 (.A1(Nb[7]), .A2(Na[20]), .ZN(n_187));
   NAND2_X1 i_188 (.A1(Nb[7]), .A2(Na[21]), .ZN(n_188));
   NAND2_X1 i_189 (.A1(Nb[7]), .A2(Na[22]), .ZN(n_189));
   NAND2_X1 i_190 (.A1(Nb[7]), .A2(Na[23]), .ZN(n_190));
   NAND2_X1 i_191 (.A1(Nb[8]), .A2(Na[0]), .ZN(n_191));
   NAND2_X1 i_192 (.A1(Nb[8]), .A2(Na[1]), .ZN(n_192));
   NAND2_X1 i_193 (.A1(Nb[8]), .A2(Na[2]), .ZN(n_193));
   NAND2_X1 i_194 (.A1(Nb[8]), .A2(Na[3]), .ZN(n_194));
   NAND2_X1 i_195 (.A1(Nb[8]), .A2(Na[4]), .ZN(n_195));
   NAND2_X1 i_196 (.A1(Nb[8]), .A2(Na[5]), .ZN(n_196));
   NAND2_X1 i_197 (.A1(Nb[8]), .A2(Na[6]), .ZN(n_197));
   NAND2_X1 i_198 (.A1(Nb[8]), .A2(Na[7]), .ZN(n_198));
   NAND2_X1 i_199 (.A1(Nb[8]), .A2(Na[8]), .ZN(n_199));
   NAND2_X1 i_200 (.A1(Nb[8]), .A2(Na[9]), .ZN(n_200));
   NAND2_X1 i_201 (.A1(Nb[8]), .A2(Na[10]), .ZN(n_201));
   NAND2_X1 i_202 (.A1(Nb[8]), .A2(Na[11]), .ZN(n_202));
   NAND2_X1 i_203 (.A1(Nb[8]), .A2(Na[12]), .ZN(n_203));
   NAND2_X1 i_204 (.A1(Nb[8]), .A2(Na[13]), .ZN(n_204));
   NAND2_X1 i_205 (.A1(Nb[8]), .A2(Na[14]), .ZN(n_205));
   NAND2_X1 i_206 (.A1(Nb[8]), .A2(Na[15]), .ZN(n_206));
   NAND2_X1 i_207 (.A1(Nb[8]), .A2(Na[16]), .ZN(n_207));
   NAND2_X1 i_208 (.A1(Nb[8]), .A2(Na[17]), .ZN(n_208));
   NAND2_X1 i_209 (.A1(Nb[8]), .A2(Na[18]), .ZN(n_209));
   NAND2_X1 i_210 (.A1(Nb[8]), .A2(Na[19]), .ZN(n_210));
   NAND2_X1 i_211 (.A1(Nb[8]), .A2(Na[20]), .ZN(n_211));
   NAND2_X1 i_212 (.A1(Nb[8]), .A2(Na[21]), .ZN(n_212));
   NAND2_X1 i_213 (.A1(Nb[8]), .A2(Na[22]), .ZN(n_213));
   NAND2_X1 i_214 (.A1(Nb[8]), .A2(Na[23]), .ZN(n_214));
   NAND2_X1 i_215 (.A1(Nb[9]), .A2(Na[0]), .ZN(n_215));
   NAND2_X1 i_216 (.A1(Nb[9]), .A2(Na[1]), .ZN(n_216));
   NAND2_X1 i_217 (.A1(Nb[9]), .A2(Na[2]), .ZN(n_217));
   NAND2_X1 i_218 (.A1(Nb[9]), .A2(Na[3]), .ZN(n_218));
   NAND2_X1 i_219 (.A1(Nb[9]), .A2(Na[4]), .ZN(n_219));
   NAND2_X1 i_220 (.A1(Nb[9]), .A2(Na[5]), .ZN(n_220));
   NAND2_X1 i_221 (.A1(Nb[9]), .A2(Na[6]), .ZN(n_221));
   NAND2_X1 i_222 (.A1(Nb[9]), .A2(Na[7]), .ZN(n_222));
   NAND2_X1 i_223 (.A1(Nb[9]), .A2(Na[8]), .ZN(n_223));
   NAND2_X1 i_224 (.A1(Nb[9]), .A2(Na[9]), .ZN(n_224));
   NAND2_X1 i_225 (.A1(Nb[9]), .A2(Na[10]), .ZN(n_225));
   NAND2_X1 i_226 (.A1(Nb[9]), .A2(Na[11]), .ZN(n_226));
   NAND2_X1 i_227 (.A1(Nb[9]), .A2(Na[12]), .ZN(n_227));
   NAND2_X1 i_228 (.A1(Nb[9]), .A2(Na[13]), .ZN(n_228));
   NAND2_X1 i_229 (.A1(Nb[9]), .A2(Na[14]), .ZN(n_229));
   NAND2_X1 i_230 (.A1(Nb[9]), .A2(Na[15]), .ZN(n_230));
   NAND2_X1 i_231 (.A1(Nb[9]), .A2(Na[16]), .ZN(n_231));
   NAND2_X1 i_232 (.A1(Nb[9]), .A2(Na[17]), .ZN(n_232));
   NAND2_X1 i_233 (.A1(Nb[9]), .A2(Na[18]), .ZN(n_233));
   NAND2_X1 i_234 (.A1(Nb[9]), .A2(Na[19]), .ZN(n_234));
   NAND2_X1 i_235 (.A1(Nb[9]), .A2(Na[20]), .ZN(n_235));
   NAND2_X1 i_236 (.A1(Nb[9]), .A2(Na[21]), .ZN(n_236));
   NAND2_X1 i_237 (.A1(Nb[9]), .A2(Na[22]), .ZN(n_237));
   NAND2_X1 i_238 (.A1(Nb[9]), .A2(Na[23]), .ZN(n_238));
   NAND2_X1 i_239 (.A1(Nb[10]), .A2(Na[0]), .ZN(n_239));
   NAND2_X1 i_240 (.A1(Nb[10]), .A2(Na[1]), .ZN(n_240));
   NAND2_X1 i_241 (.A1(Nb[10]), .A2(Na[2]), .ZN(n_241));
   NAND2_X1 i_242 (.A1(Nb[10]), .A2(Na[3]), .ZN(n_242));
   NAND2_X1 i_243 (.A1(Nb[10]), .A2(Na[4]), .ZN(n_243));
   NAND2_X1 i_244 (.A1(Nb[10]), .A2(Na[5]), .ZN(n_244));
   NAND2_X1 i_245 (.A1(Nb[10]), .A2(Na[6]), .ZN(n_245));
   NAND2_X1 i_246 (.A1(Nb[10]), .A2(Na[7]), .ZN(n_246));
   NAND2_X1 i_247 (.A1(Nb[10]), .A2(Na[8]), .ZN(n_247));
   NAND2_X1 i_248 (.A1(Nb[10]), .A2(Na[9]), .ZN(n_248));
   NAND2_X1 i_249 (.A1(Nb[10]), .A2(Na[10]), .ZN(n_249));
   NAND2_X1 i_250 (.A1(Nb[10]), .A2(Na[11]), .ZN(n_250));
   NAND2_X1 i_251 (.A1(Nb[10]), .A2(Na[12]), .ZN(n_251));
   NAND2_X1 i_252 (.A1(Nb[10]), .A2(Na[13]), .ZN(n_252));
   NAND2_X1 i_253 (.A1(Nb[10]), .A2(Na[14]), .ZN(n_253));
   NAND2_X1 i_254 (.A1(Nb[10]), .A2(Na[15]), .ZN(n_254));
   NAND2_X1 i_255 (.A1(Nb[10]), .A2(Na[16]), .ZN(n_255));
   NAND2_X1 i_256 (.A1(Nb[10]), .A2(Na[17]), .ZN(n_256));
   NAND2_X1 i_257 (.A1(Nb[10]), .A2(Na[18]), .ZN(n_257));
   NAND2_X1 i_258 (.A1(Nb[10]), .A2(Na[19]), .ZN(n_258));
   NAND2_X1 i_259 (.A1(Nb[10]), .A2(Na[20]), .ZN(n_259));
   NAND2_X1 i_260 (.A1(Nb[10]), .A2(Na[21]), .ZN(n_260));
   NAND2_X1 i_261 (.A1(Nb[10]), .A2(Na[22]), .ZN(n_261));
   NAND2_X1 i_262 (.A1(Nb[10]), .A2(Na[23]), .ZN(n_262));
   NAND2_X1 i_263 (.A1(Nb[11]), .A2(Na[0]), .ZN(n_263));
   NAND2_X1 i_264 (.A1(Nb[11]), .A2(Na[1]), .ZN(n_264));
   NAND2_X1 i_265 (.A1(Nb[11]), .A2(Na[2]), .ZN(n_265));
   NAND2_X1 i_266 (.A1(Nb[11]), .A2(Na[3]), .ZN(n_266));
   NAND2_X1 i_267 (.A1(Nb[11]), .A2(Na[4]), .ZN(n_267));
   NAND2_X1 i_268 (.A1(Nb[11]), .A2(Na[5]), .ZN(n_268));
   NAND2_X1 i_269 (.A1(Nb[11]), .A2(Na[6]), .ZN(n_269));
   NAND2_X1 i_270 (.A1(Nb[11]), .A2(Na[7]), .ZN(n_270));
   NAND2_X1 i_271 (.A1(Nb[11]), .A2(Na[8]), .ZN(n_271));
   NAND2_X1 i_272 (.A1(Nb[11]), .A2(Na[9]), .ZN(n_272));
   NAND2_X1 i_273 (.A1(Nb[11]), .A2(Na[10]), .ZN(n_273));
   NAND2_X1 i_274 (.A1(Nb[11]), .A2(Na[11]), .ZN(n_274));
   NAND2_X1 i_275 (.A1(Nb[11]), .A2(Na[12]), .ZN(n_275));
   NAND2_X1 i_276 (.A1(Nb[11]), .A2(Na[13]), .ZN(n_276));
   NAND2_X1 i_277 (.A1(Nb[11]), .A2(Na[14]), .ZN(n_277));
   NAND2_X1 i_278 (.A1(Nb[11]), .A2(Na[15]), .ZN(n_278));
   NAND2_X1 i_279 (.A1(Nb[11]), .A2(Na[16]), .ZN(n_279));
   NAND2_X1 i_280 (.A1(Nb[11]), .A2(Na[17]), .ZN(n_280));
   NAND2_X1 i_281 (.A1(Nb[11]), .A2(Na[18]), .ZN(n_281));
   NAND2_X1 i_282 (.A1(Nb[11]), .A2(Na[19]), .ZN(n_282));
   NAND2_X1 i_283 (.A1(Nb[11]), .A2(Na[20]), .ZN(n_283));
   NAND2_X1 i_284 (.A1(Nb[11]), .A2(Na[21]), .ZN(n_284));
   NAND2_X1 i_285 (.A1(Nb[11]), .A2(Na[22]), .ZN(n_285));
   NAND2_X1 i_286 (.A1(Nb[11]), .A2(Na[23]), .ZN(n_286));
   NAND2_X1 i_287 (.A1(Nb[12]), .A2(Na[0]), .ZN(n_287));
   NAND2_X1 i_288 (.A1(Nb[12]), .A2(Na[1]), .ZN(n_288));
   NAND2_X1 i_289 (.A1(Nb[12]), .A2(Na[2]), .ZN(n_289));
   NAND2_X1 i_290 (.A1(Nb[12]), .A2(Na[3]), .ZN(n_290));
   NAND2_X1 i_291 (.A1(Nb[12]), .A2(Na[4]), .ZN(n_291));
   NAND2_X1 i_292 (.A1(Nb[12]), .A2(Na[5]), .ZN(n_292));
   NAND2_X1 i_293 (.A1(Nb[12]), .A2(Na[6]), .ZN(n_293));
   NAND2_X1 i_294 (.A1(Nb[12]), .A2(Na[7]), .ZN(n_294));
   NAND2_X1 i_295 (.A1(Nb[12]), .A2(Na[8]), .ZN(n_295));
   NAND2_X1 i_296 (.A1(Nb[12]), .A2(Na[9]), .ZN(n_296));
   NAND2_X1 i_297 (.A1(Nb[12]), .A2(Na[10]), .ZN(n_297));
   NAND2_X1 i_298 (.A1(Nb[12]), .A2(Na[11]), .ZN(n_298));
   NAND2_X1 i_299 (.A1(Nb[12]), .A2(Na[12]), .ZN(n_299));
   NAND2_X1 i_300 (.A1(Nb[12]), .A2(Na[13]), .ZN(n_300));
   NAND2_X1 i_301 (.A1(Nb[12]), .A2(Na[14]), .ZN(n_301));
   NAND2_X1 i_302 (.A1(Nb[12]), .A2(Na[15]), .ZN(n_302));
   NAND2_X1 i_303 (.A1(Nb[12]), .A2(Na[16]), .ZN(n_303));
   NAND2_X1 i_304 (.A1(Nb[12]), .A2(Na[17]), .ZN(n_304));
   NAND2_X1 i_305 (.A1(Nb[12]), .A2(Na[18]), .ZN(n_305));
   NAND2_X1 i_306 (.A1(Nb[12]), .A2(Na[19]), .ZN(n_306));
   NAND2_X1 i_307 (.A1(Nb[12]), .A2(Na[20]), .ZN(n_307));
   NAND2_X1 i_308 (.A1(Nb[12]), .A2(Na[21]), .ZN(n_308));
   NAND2_X1 i_309 (.A1(Nb[12]), .A2(Na[22]), .ZN(n_309));
   NAND2_X1 i_310 (.A1(Nb[12]), .A2(Na[23]), .ZN(n_310));
   NAND2_X1 i_311 (.A1(Nb[13]), .A2(Na[0]), .ZN(n_311));
   NAND2_X1 i_312 (.A1(Nb[13]), .A2(Na[1]), .ZN(n_312));
   NAND2_X1 i_313 (.A1(Nb[13]), .A2(Na[2]), .ZN(n_313));
   NAND2_X1 i_314 (.A1(Nb[13]), .A2(Na[3]), .ZN(n_314));
   NAND2_X1 i_315 (.A1(Nb[13]), .A2(Na[4]), .ZN(n_315));
   NAND2_X1 i_316 (.A1(Nb[13]), .A2(Na[5]), .ZN(n_316));
   NAND2_X1 i_317 (.A1(Nb[13]), .A2(Na[6]), .ZN(n_317));
   NAND2_X1 i_318 (.A1(Nb[13]), .A2(Na[7]), .ZN(n_318));
   NAND2_X1 i_319 (.A1(Nb[13]), .A2(Na[8]), .ZN(n_319));
   NAND2_X1 i_320 (.A1(Nb[13]), .A2(Na[9]), .ZN(n_320));
   NAND2_X1 i_321 (.A1(Nb[13]), .A2(Na[10]), .ZN(n_321));
   NAND2_X1 i_322 (.A1(Nb[13]), .A2(Na[11]), .ZN(n_322));
   NAND2_X1 i_323 (.A1(Nb[13]), .A2(Na[12]), .ZN(n_323));
   NAND2_X1 i_324 (.A1(Nb[13]), .A2(Na[13]), .ZN(n_324));
   NAND2_X1 i_325 (.A1(Nb[13]), .A2(Na[14]), .ZN(n_325));
   NAND2_X1 i_326 (.A1(Nb[13]), .A2(Na[15]), .ZN(n_326));
   NAND2_X1 i_327 (.A1(Nb[13]), .A2(Na[16]), .ZN(n_327));
   NAND2_X1 i_328 (.A1(Nb[13]), .A2(Na[17]), .ZN(n_328));
   NAND2_X1 i_329 (.A1(Nb[13]), .A2(Na[18]), .ZN(n_329));
   NAND2_X1 i_330 (.A1(Nb[13]), .A2(Na[19]), .ZN(n_330));
   NAND2_X1 i_331 (.A1(Nb[13]), .A2(Na[20]), .ZN(n_331));
   NAND2_X1 i_332 (.A1(Nb[13]), .A2(Na[21]), .ZN(n_332));
   NAND2_X1 i_333 (.A1(Nb[13]), .A2(Na[22]), .ZN(n_333));
   NAND2_X1 i_334 (.A1(Nb[13]), .A2(Na[23]), .ZN(n_334));
   NAND2_X1 i_335 (.A1(Nb[14]), .A2(Na[0]), .ZN(n_335));
   NAND2_X1 i_336 (.A1(Nb[14]), .A2(Na[1]), .ZN(n_336));
   NAND2_X1 i_337 (.A1(Nb[14]), .A2(Na[2]), .ZN(n_337));
   NAND2_X1 i_338 (.A1(Nb[14]), .A2(Na[3]), .ZN(n_338));
   NAND2_X1 i_339 (.A1(Nb[14]), .A2(Na[4]), .ZN(n_339));
   NAND2_X1 i_340 (.A1(Nb[14]), .A2(Na[5]), .ZN(n_340));
   NAND2_X1 i_341 (.A1(Nb[14]), .A2(Na[6]), .ZN(n_341));
   NAND2_X1 i_342 (.A1(Nb[14]), .A2(Na[7]), .ZN(n_342));
   NAND2_X1 i_343 (.A1(Nb[14]), .A2(Na[8]), .ZN(n_343));
   NAND2_X1 i_344 (.A1(Nb[14]), .A2(Na[9]), .ZN(n_344));
   NAND2_X1 i_345 (.A1(Nb[14]), .A2(Na[10]), .ZN(n_345));
   NAND2_X1 i_346 (.A1(Nb[14]), .A2(Na[11]), .ZN(n_346));
   NAND2_X1 i_347 (.A1(Nb[14]), .A2(Na[12]), .ZN(n_347));
   NAND2_X1 i_348 (.A1(Nb[14]), .A2(Na[13]), .ZN(n_348));
   NAND2_X1 i_349 (.A1(Nb[14]), .A2(Na[14]), .ZN(n_349));
   NAND2_X1 i_350 (.A1(Nb[14]), .A2(Na[15]), .ZN(n_350));
   NAND2_X1 i_351 (.A1(Nb[14]), .A2(Na[16]), .ZN(n_351));
   NAND2_X1 i_352 (.A1(Nb[14]), .A2(Na[17]), .ZN(n_352));
   NAND2_X1 i_353 (.A1(Nb[14]), .A2(Na[18]), .ZN(n_353));
   NAND2_X1 i_354 (.A1(Nb[14]), .A2(Na[19]), .ZN(n_354));
   NAND2_X1 i_355 (.A1(Nb[14]), .A2(Na[20]), .ZN(n_355));
   NAND2_X1 i_356 (.A1(Nb[14]), .A2(Na[21]), .ZN(n_356));
   NAND2_X1 i_357 (.A1(Nb[14]), .A2(Na[22]), .ZN(n_357));
   NAND2_X1 i_358 (.A1(Nb[14]), .A2(Na[23]), .ZN(n_358));
   NAND2_X1 i_359 (.A1(Nb[15]), .A2(Na[0]), .ZN(n_359));
   NAND2_X1 i_360 (.A1(Nb[15]), .A2(Na[1]), .ZN(n_360));
   NAND2_X1 i_361 (.A1(Nb[15]), .A2(Na[2]), .ZN(n_361));
   NAND2_X1 i_362 (.A1(Nb[15]), .A2(Na[3]), .ZN(n_362));
   NAND2_X1 i_363 (.A1(Nb[15]), .A2(Na[4]), .ZN(n_363));
   NAND2_X1 i_364 (.A1(Nb[15]), .A2(Na[5]), .ZN(n_364));
   NAND2_X1 i_365 (.A1(Nb[15]), .A2(Na[6]), .ZN(n_365));
   NAND2_X1 i_366 (.A1(Nb[15]), .A2(Na[7]), .ZN(n_366));
   NAND2_X1 i_367 (.A1(Nb[15]), .A2(Na[8]), .ZN(n_367));
   NAND2_X1 i_368 (.A1(Nb[15]), .A2(Na[9]), .ZN(n_368));
   NAND2_X1 i_369 (.A1(Nb[15]), .A2(Na[10]), .ZN(n_369));
   NAND2_X1 i_370 (.A1(Nb[15]), .A2(Na[11]), .ZN(n_370));
   NAND2_X1 i_371 (.A1(Nb[15]), .A2(Na[12]), .ZN(n_371));
   NAND2_X1 i_372 (.A1(Nb[15]), .A2(Na[13]), .ZN(n_372));
   NAND2_X1 i_373 (.A1(Nb[15]), .A2(Na[14]), .ZN(n_373));
   NAND2_X1 i_374 (.A1(Nb[15]), .A2(Na[15]), .ZN(n_374));
   NAND2_X1 i_375 (.A1(Nb[15]), .A2(Na[16]), .ZN(n_375));
   NAND2_X1 i_376 (.A1(Nb[15]), .A2(Na[17]), .ZN(n_376));
   NAND2_X1 i_377 (.A1(Nb[15]), .A2(Na[18]), .ZN(n_377));
   NAND2_X1 i_378 (.A1(Nb[15]), .A2(Na[19]), .ZN(n_378));
   NAND2_X1 i_379 (.A1(Nb[15]), .A2(Na[20]), .ZN(n_379));
   NAND2_X1 i_380 (.A1(Nb[15]), .A2(Na[21]), .ZN(n_380));
   NAND2_X1 i_381 (.A1(Nb[15]), .A2(Na[22]), .ZN(n_381));
   NAND2_X1 i_382 (.A1(Nb[15]), .A2(Na[23]), .ZN(n_382));
   NAND2_X1 i_383 (.A1(Nb[16]), .A2(Na[0]), .ZN(n_383));
   NAND2_X1 i_384 (.A1(Nb[16]), .A2(Na[1]), .ZN(n_384));
   NAND2_X1 i_385 (.A1(Nb[16]), .A2(Na[2]), .ZN(n_385));
   NAND2_X1 i_386 (.A1(Nb[16]), .A2(Na[3]), .ZN(n_386));
   NAND2_X1 i_387 (.A1(Nb[16]), .A2(Na[4]), .ZN(n_387));
   NAND2_X1 i_388 (.A1(Nb[16]), .A2(Na[5]), .ZN(n_388));
   NAND2_X1 i_389 (.A1(Nb[16]), .A2(Na[6]), .ZN(n_389));
   NAND2_X1 i_390 (.A1(Nb[16]), .A2(Na[7]), .ZN(n_390));
   NAND2_X1 i_391 (.A1(Nb[16]), .A2(Na[8]), .ZN(n_391));
   NAND2_X1 i_392 (.A1(Nb[16]), .A2(Na[9]), .ZN(n_392));
   NAND2_X1 i_393 (.A1(Nb[16]), .A2(Na[10]), .ZN(n_393));
   NAND2_X1 i_394 (.A1(Nb[16]), .A2(Na[11]), .ZN(n_394));
   NAND2_X1 i_395 (.A1(Nb[16]), .A2(Na[12]), .ZN(n_395));
   NAND2_X1 i_396 (.A1(Nb[16]), .A2(Na[13]), .ZN(n_396));
   NAND2_X1 i_397 (.A1(Nb[16]), .A2(Na[14]), .ZN(n_397));
   NAND2_X1 i_398 (.A1(Nb[16]), .A2(Na[15]), .ZN(n_398));
   NAND2_X1 i_399 (.A1(Nb[16]), .A2(Na[16]), .ZN(n_399));
   NAND2_X1 i_400 (.A1(Nb[16]), .A2(Na[17]), .ZN(n_400));
   NAND2_X1 i_401 (.A1(Nb[16]), .A2(Na[18]), .ZN(n_401));
   NAND2_X1 i_402 (.A1(Nb[16]), .A2(Na[19]), .ZN(n_402));
   NAND2_X1 i_403 (.A1(Nb[16]), .A2(Na[20]), .ZN(n_403));
   NAND2_X1 i_404 (.A1(Nb[16]), .A2(Na[21]), .ZN(n_404));
   NAND2_X1 i_405 (.A1(Nb[16]), .A2(Na[22]), .ZN(n_405));
   NAND2_X1 i_406 (.A1(Nb[16]), .A2(Na[23]), .ZN(n_406));
   NAND2_X1 i_407 (.A1(Nb[17]), .A2(Na[0]), .ZN(n_407));
   NAND2_X1 i_408 (.A1(Nb[17]), .A2(Na[1]), .ZN(n_408));
   NAND2_X1 i_409 (.A1(Nb[17]), .A2(Na[2]), .ZN(n_409));
   NAND2_X1 i_410 (.A1(Nb[17]), .A2(Na[3]), .ZN(n_410));
   NAND2_X1 i_411 (.A1(Nb[17]), .A2(Na[4]), .ZN(n_411));
   NAND2_X1 i_412 (.A1(Nb[17]), .A2(Na[5]), .ZN(n_412));
   NAND2_X1 i_413 (.A1(Nb[17]), .A2(Na[6]), .ZN(n_413));
   NAND2_X1 i_414 (.A1(Nb[17]), .A2(Na[7]), .ZN(n_414));
   NAND2_X1 i_415 (.A1(Nb[17]), .A2(Na[8]), .ZN(n_415));
   NAND2_X1 i_416 (.A1(Nb[17]), .A2(Na[9]), .ZN(n_416));
   NAND2_X1 i_417 (.A1(Nb[17]), .A2(Na[10]), .ZN(n_417));
   NAND2_X1 i_418 (.A1(Nb[17]), .A2(Na[11]), .ZN(n_418));
   NAND2_X1 i_419 (.A1(Nb[17]), .A2(Na[12]), .ZN(n_419));
   NAND2_X1 i_420 (.A1(Nb[17]), .A2(Na[13]), .ZN(n_420));
   NAND2_X1 i_421 (.A1(Nb[17]), .A2(Na[14]), .ZN(n_421));
   NAND2_X1 i_422 (.A1(Nb[17]), .A2(Na[15]), .ZN(n_422));
   NAND2_X1 i_423 (.A1(Nb[17]), .A2(Na[16]), .ZN(n_423));
   NAND2_X1 i_424 (.A1(Nb[17]), .A2(Na[17]), .ZN(n_424));
   NAND2_X1 i_425 (.A1(Nb[17]), .A2(Na[18]), .ZN(n_425));
   NAND2_X1 i_426 (.A1(Nb[17]), .A2(Na[19]), .ZN(n_426));
   NAND2_X1 i_427 (.A1(Nb[17]), .A2(Na[20]), .ZN(n_427));
   NAND2_X1 i_428 (.A1(Nb[17]), .A2(Na[21]), .ZN(n_428));
   NAND2_X1 i_429 (.A1(Nb[17]), .A2(Na[22]), .ZN(n_429));
   NAND2_X1 i_430 (.A1(Nb[17]), .A2(Na[23]), .ZN(n_430));
   NAND2_X1 i_431 (.A1(Nb[18]), .A2(Na[0]), .ZN(n_431));
   NAND2_X1 i_432 (.A1(Nb[18]), .A2(Na[1]), .ZN(n_432));
   NAND2_X1 i_433 (.A1(Nb[18]), .A2(Na[2]), .ZN(n_433));
   NAND2_X1 i_434 (.A1(Nb[18]), .A2(Na[3]), .ZN(n_434));
   NAND2_X1 i_435 (.A1(Nb[18]), .A2(Na[4]), .ZN(n_435));
   NAND2_X1 i_436 (.A1(Nb[18]), .A2(Na[5]), .ZN(n_436));
   NAND2_X1 i_437 (.A1(Nb[18]), .A2(Na[6]), .ZN(n_437));
   NAND2_X1 i_438 (.A1(Nb[18]), .A2(Na[7]), .ZN(n_438));
   NAND2_X1 i_439 (.A1(Nb[18]), .A2(Na[8]), .ZN(n_439));
   NAND2_X1 i_440 (.A1(Nb[18]), .A2(Na[9]), .ZN(n_440));
   NAND2_X1 i_441 (.A1(Nb[18]), .A2(Na[10]), .ZN(n_441));
   NAND2_X1 i_442 (.A1(Nb[18]), .A2(Na[11]), .ZN(n_442));
   NAND2_X1 i_443 (.A1(Nb[18]), .A2(Na[12]), .ZN(n_443));
   NAND2_X1 i_444 (.A1(Nb[18]), .A2(Na[13]), .ZN(n_444));
   NAND2_X1 i_445 (.A1(Nb[18]), .A2(Na[14]), .ZN(n_445));
   NAND2_X1 i_446 (.A1(Nb[18]), .A2(Na[15]), .ZN(n_446));
   NAND2_X1 i_447 (.A1(Nb[18]), .A2(Na[16]), .ZN(n_447));
   NAND2_X1 i_448 (.A1(Nb[18]), .A2(Na[17]), .ZN(n_448));
   NAND2_X1 i_449 (.A1(Nb[18]), .A2(Na[18]), .ZN(n_449));
   NAND2_X1 i_450 (.A1(Nb[18]), .A2(Na[19]), .ZN(n_450));
   NAND2_X1 i_451 (.A1(Nb[18]), .A2(Na[20]), .ZN(n_451));
   NAND2_X1 i_452 (.A1(Nb[18]), .A2(Na[21]), .ZN(n_452));
   NAND2_X1 i_453 (.A1(Nb[18]), .A2(Na[22]), .ZN(n_453));
   NAND2_X1 i_454 (.A1(Nb[18]), .A2(Na[23]), .ZN(n_454));
   NAND2_X1 i_455 (.A1(Nb[19]), .A2(Na[0]), .ZN(n_455));
   NAND2_X1 i_456 (.A1(Nb[19]), .A2(Na[1]), .ZN(n_456));
   NAND2_X1 i_457 (.A1(Nb[19]), .A2(Na[2]), .ZN(n_457));
   NAND2_X1 i_458 (.A1(Nb[19]), .A2(Na[3]), .ZN(n_458));
   NAND2_X1 i_459 (.A1(Nb[19]), .A2(Na[4]), .ZN(n_459));
   NAND2_X1 i_460 (.A1(Nb[19]), .A2(Na[5]), .ZN(n_460));
   NAND2_X1 i_461 (.A1(Nb[19]), .A2(Na[6]), .ZN(n_461));
   NAND2_X1 i_462 (.A1(Nb[19]), .A2(Na[7]), .ZN(n_462));
   NAND2_X1 i_463 (.A1(Nb[19]), .A2(Na[8]), .ZN(n_463));
   NAND2_X1 i_464 (.A1(Nb[19]), .A2(Na[9]), .ZN(n_464));
   NAND2_X1 i_465 (.A1(Nb[19]), .A2(Na[10]), .ZN(n_465));
   NAND2_X1 i_466 (.A1(Nb[19]), .A2(Na[11]), .ZN(n_466));
   NAND2_X1 i_467 (.A1(Nb[19]), .A2(Na[12]), .ZN(n_467));
   NAND2_X1 i_468 (.A1(Nb[19]), .A2(Na[13]), .ZN(n_468));
   NAND2_X1 i_469 (.A1(Nb[19]), .A2(Na[14]), .ZN(n_469));
   NAND2_X1 i_470 (.A1(Nb[19]), .A2(Na[15]), .ZN(n_470));
   NAND2_X1 i_471 (.A1(Nb[19]), .A2(Na[16]), .ZN(n_471));
   NAND2_X1 i_472 (.A1(Nb[19]), .A2(Na[17]), .ZN(n_472));
   NAND2_X1 i_473 (.A1(Nb[19]), .A2(Na[18]), .ZN(n_473));
   NAND2_X1 i_474 (.A1(Nb[19]), .A2(Na[19]), .ZN(n_474));
   NAND2_X1 i_475 (.A1(Nb[19]), .A2(Na[20]), .ZN(n_475));
   NAND2_X1 i_476 (.A1(Nb[19]), .A2(Na[21]), .ZN(n_476));
   NAND2_X1 i_477 (.A1(Nb[19]), .A2(Na[22]), .ZN(n_477));
   NAND2_X1 i_478 (.A1(Nb[19]), .A2(Na[23]), .ZN(n_478));
   NAND2_X1 i_479 (.A1(Nb[20]), .A2(Na[0]), .ZN(n_479));
   NAND2_X1 i_480 (.A1(Nb[20]), .A2(Na[1]), .ZN(n_480));
   NAND2_X1 i_481 (.A1(Nb[20]), .A2(Na[2]), .ZN(n_481));
   NAND2_X1 i_482 (.A1(Nb[20]), .A2(Na[3]), .ZN(n_482));
   NAND2_X1 i_483 (.A1(Nb[20]), .A2(Na[4]), .ZN(n_483));
   NAND2_X1 i_484 (.A1(Nb[20]), .A2(Na[5]), .ZN(n_484));
   NAND2_X1 i_485 (.A1(Nb[20]), .A2(Na[6]), .ZN(n_485));
   NAND2_X1 i_486 (.A1(Nb[20]), .A2(Na[7]), .ZN(n_486));
   NAND2_X1 i_487 (.A1(Nb[20]), .A2(Na[8]), .ZN(n_487));
   NAND2_X1 i_488 (.A1(Nb[20]), .A2(Na[9]), .ZN(n_488));
   NAND2_X1 i_489 (.A1(Nb[20]), .A2(Na[10]), .ZN(n_489));
   NAND2_X1 i_490 (.A1(Nb[20]), .A2(Na[11]), .ZN(n_490));
   NAND2_X1 i_491 (.A1(Nb[20]), .A2(Na[12]), .ZN(n_491));
   NAND2_X1 i_492 (.A1(Nb[20]), .A2(Na[13]), .ZN(n_492));
   NAND2_X1 i_493 (.A1(Nb[20]), .A2(Na[14]), .ZN(n_493));
   NAND2_X1 i_494 (.A1(Nb[20]), .A2(Na[15]), .ZN(n_494));
   NAND2_X1 i_495 (.A1(Nb[20]), .A2(Na[16]), .ZN(n_495));
   NAND2_X1 i_496 (.A1(Nb[20]), .A2(Na[17]), .ZN(n_496));
   NAND2_X1 i_497 (.A1(Nb[20]), .A2(Na[18]), .ZN(n_497));
   NAND2_X1 i_498 (.A1(Nb[20]), .A2(Na[19]), .ZN(n_498));
   NAND2_X1 i_499 (.A1(Nb[20]), .A2(Na[20]), .ZN(n_499));
   NAND2_X1 i_500 (.A1(Nb[20]), .A2(Na[21]), .ZN(n_500));
   NAND2_X1 i_501 (.A1(Nb[20]), .A2(Na[22]), .ZN(n_501));
   NAND2_X1 i_502 (.A1(Nb[20]), .A2(Na[23]), .ZN(n_502));
   NAND2_X1 i_503 (.A1(Nb[21]), .A2(Na[0]), .ZN(n_503));
   NAND2_X1 i_504 (.A1(Nb[21]), .A2(Na[1]), .ZN(n_504));
   NAND2_X1 i_505 (.A1(Nb[21]), .A2(Na[2]), .ZN(n_505));
   NAND2_X1 i_506 (.A1(Nb[21]), .A2(Na[3]), .ZN(n_506));
   NAND2_X1 i_507 (.A1(Nb[21]), .A2(Na[4]), .ZN(n_507));
   NAND2_X1 i_508 (.A1(Nb[21]), .A2(Na[5]), .ZN(n_508));
   NAND2_X1 i_509 (.A1(Nb[21]), .A2(Na[6]), .ZN(n_509));
   NAND2_X1 i_510 (.A1(Nb[21]), .A2(Na[7]), .ZN(n_510));
   NAND2_X1 i_511 (.A1(Nb[21]), .A2(Na[8]), .ZN(n_511));
   NAND2_X1 i_512 (.A1(Nb[21]), .A2(Na[9]), .ZN(n_512));
   NAND2_X1 i_513 (.A1(Nb[21]), .A2(Na[10]), .ZN(n_513));
   NAND2_X1 i_514 (.A1(Nb[21]), .A2(Na[11]), .ZN(n_514));
   NAND2_X1 i_515 (.A1(Nb[21]), .A2(Na[12]), .ZN(n_515));
   NAND2_X1 i_516 (.A1(Nb[21]), .A2(Na[13]), .ZN(n_516));
   NAND2_X1 i_517 (.A1(Nb[21]), .A2(Na[14]), .ZN(n_517));
   NAND2_X1 i_518 (.A1(Nb[21]), .A2(Na[15]), .ZN(n_518));
   NAND2_X1 i_519 (.A1(Nb[21]), .A2(Na[16]), .ZN(n_519));
   NAND2_X1 i_520 (.A1(Nb[21]), .A2(Na[17]), .ZN(n_520));
   NAND2_X1 i_521 (.A1(Nb[21]), .A2(Na[18]), .ZN(n_521));
   NAND2_X1 i_522 (.A1(Nb[21]), .A2(Na[19]), .ZN(n_522));
   NAND2_X1 i_523 (.A1(Nb[21]), .A2(Na[20]), .ZN(n_523));
   NAND2_X1 i_524 (.A1(Nb[21]), .A2(Na[21]), .ZN(n_524));
   NAND2_X1 i_525 (.A1(Nb[21]), .A2(Na[22]), .ZN(n_525));
   NAND2_X1 i_526 (.A1(Nb[21]), .A2(Na[23]), .ZN(n_526));
   NAND2_X1 i_527 (.A1(Nb[22]), .A2(Na[0]), .ZN(n_527));
   NAND2_X1 i_528 (.A1(Nb[22]), .A2(Na[1]), .ZN(n_528));
   NAND2_X1 i_529 (.A1(Nb[22]), .A2(Na[2]), .ZN(n_529));
   NAND2_X1 i_530 (.A1(Nb[22]), .A2(Na[3]), .ZN(n_530));
   NAND2_X1 i_531 (.A1(Nb[22]), .A2(Na[4]), .ZN(n_531));
   NAND2_X1 i_532 (.A1(Nb[22]), .A2(Na[5]), .ZN(n_532));
   NAND2_X1 i_533 (.A1(Nb[22]), .A2(Na[6]), .ZN(n_533));
   NAND2_X1 i_534 (.A1(Nb[22]), .A2(Na[7]), .ZN(n_534));
   NAND2_X1 i_535 (.A1(Nb[22]), .A2(Na[8]), .ZN(n_535));
   NAND2_X1 i_536 (.A1(Nb[22]), .A2(Na[9]), .ZN(n_536));
   NAND2_X1 i_537 (.A1(Nb[22]), .A2(Na[10]), .ZN(n_537));
   NAND2_X1 i_538 (.A1(Nb[22]), .A2(Na[11]), .ZN(n_538));
   NAND2_X1 i_539 (.A1(Nb[22]), .A2(Na[12]), .ZN(n_539));
   NAND2_X1 i_540 (.A1(Nb[22]), .A2(Na[13]), .ZN(n_540));
   NAND2_X1 i_541 (.A1(Nb[22]), .A2(Na[14]), .ZN(n_541));
   NAND2_X1 i_542 (.A1(Nb[22]), .A2(Na[15]), .ZN(n_542));
   NAND2_X1 i_543 (.A1(Nb[22]), .A2(Na[16]), .ZN(n_543));
   NAND2_X1 i_544 (.A1(Nb[22]), .A2(Na[17]), .ZN(n_544));
   NAND2_X1 i_545 (.A1(Nb[22]), .A2(Na[18]), .ZN(n_545));
   NAND2_X1 i_546 (.A1(Nb[22]), .A2(Na[19]), .ZN(n_546));
   NAND2_X1 i_547 (.A1(Nb[22]), .A2(Na[20]), .ZN(n_547));
   NAND2_X1 i_548 (.A1(Nb[22]), .A2(Na[21]), .ZN(n_548));
   NAND2_X1 i_549 (.A1(Nb[22]), .A2(Na[22]), .ZN(n_549));
   NAND2_X1 i_550 (.A1(Nb[22]), .A2(Na[23]), .ZN(n_550));
   NAND2_X1 i_551 (.A1(Nb[23]), .A2(Na[0]), .ZN(n_551));
   NAND2_X1 i_552 (.A1(Nb[23]), .A2(Na[1]), .ZN(n_552));
   NAND2_X1 i_553 (.A1(Nb[23]), .A2(Na[2]), .ZN(n_553));
   NAND2_X1 i_554 (.A1(Nb[23]), .A2(Na[3]), .ZN(n_554));
   NAND2_X1 i_555 (.A1(Nb[23]), .A2(Na[4]), .ZN(n_555));
   NAND2_X1 i_556 (.A1(Nb[23]), .A2(Na[5]), .ZN(n_556));
   NAND2_X1 i_557 (.A1(Nb[23]), .A2(Na[6]), .ZN(n_557));
   NAND2_X1 i_558 (.A1(Nb[23]), .A2(Na[7]), .ZN(n_558));
   NAND2_X1 i_559 (.A1(Nb[23]), .A2(Na[8]), .ZN(n_559));
   NAND2_X1 i_560 (.A1(Nb[23]), .A2(Na[9]), .ZN(n_560));
   NAND2_X1 i_561 (.A1(Nb[23]), .A2(Na[10]), .ZN(n_561));
   NAND2_X1 i_562 (.A1(Nb[23]), .A2(Na[11]), .ZN(n_562));
   NAND2_X1 i_563 (.A1(Nb[23]), .A2(Na[12]), .ZN(n_563));
   NAND2_X1 i_564 (.A1(Nb[23]), .A2(Na[13]), .ZN(n_564));
   NAND2_X1 i_565 (.A1(Nb[23]), .A2(Na[14]), .ZN(n_565));
   NAND2_X1 i_566 (.A1(Nb[23]), .A2(Na[15]), .ZN(n_566));
   NAND2_X1 i_567 (.A1(Nb[23]), .A2(Na[16]), .ZN(n_567));
   NAND2_X1 i_568 (.A1(Nb[23]), .A2(Na[17]), .ZN(n_568));
   NAND2_X1 i_569 (.A1(Nb[23]), .A2(Na[18]), .ZN(n_569));
   NAND2_X1 i_570 (.A1(Nb[23]), .A2(Na[19]), .ZN(n_570));
   NAND2_X1 i_571 (.A1(Nb[23]), .A2(Na[20]), .ZN(n_571));
   NAND2_X1 i_572 (.A1(Nb[23]), .A2(Na[21]), .ZN(n_572));
   NAND2_X1 i_573 (.A1(Nb[23]), .A2(Na[22]), .ZN(n_573));
   NAND2_X1 i_574 (.A1(Nb[23]), .A2(Na[23]), .ZN(n_574));
   XNOR2_X1 i_575 (.A(n_47), .B(n_24), .ZN(n_575));
   INV_X1 i_576 (.A(n_575), .ZN(n_576));
   NOR2_X1 i_577 (.A1(n_24), .A2(n_47), .ZN(n_577));
   XNOR2_X1 i_578 (.A(n_71), .B(n_48), .ZN(n_578));
   XNOR2_X1 i_579 (.A(n_578), .B(n_25), .ZN(n_579));
   INV_X1 i_580 (.A(n_579), .ZN(n_580));
   OR3_X1 i_581 (.A1(n_582), .A2(n_583), .A3(n_584), .ZN(n_581));
   NOR2_X1 i_582 (.A1(n_48), .A2(n_71), .ZN(n_582));
   NOR2_X1 i_583 (.A1(n_25), .A2(n_71), .ZN(n_583));
   NOR2_X1 i_584 (.A1(n_25), .A2(n_48), .ZN(n_584));
   XNOR2_X1 i_585 (.A(n_2), .B(n_577), .ZN(n_585));
   NOR2_X1 i_586 (.A1(n_2), .A2(n_587), .ZN(n_586));
   INV_X1 i_587 (.A(n_577), .ZN(n_587));
   XNOR2_X1 i_588 (.A(n_95), .B(n_72), .ZN(n_588));
   XNOR2_X1 i_589 (.A(n_588), .B(n_49), .ZN(n_589));
   INV_X1 i_590 (.A(n_589), .ZN(n_590));
   OR3_X1 i_591 (.A1(n_592), .A2(n_593), .A3(n_594), .ZN(n_591));
   NOR2_X1 i_592 (.A1(n_72), .A2(n_95), .ZN(n_592));
   NOR2_X1 i_593 (.A1(n_49), .A2(n_95), .ZN(n_593));
   NOR2_X1 i_594 (.A1(n_49), .A2(n_72), .ZN(n_594));
   XNOR2_X1 i_595 (.A(n_26), .B(n_3), .ZN(n_595));
   XNOR2_X1 i_596 (.A(n_595), .B(n_586), .ZN(n_596));
   NAND3_X1 i_597 (.A1(n_598), .A2(n_599), .A3(n_601), .ZN(n_597));
   OR2_X1 i_598 (.A1(n_3), .A2(n_26), .ZN(n_598));
   NAND2_X1 i_599 (.A1(n_586), .A2(n_600), .ZN(n_599));
   INV_X1 i_600 (.A(n_26), .ZN(n_600));
   NAND2_X1 i_601 (.A1(n_586), .A2(n_602), .ZN(n_601));
   INV_X1 i_602 (.A(n_3), .ZN(n_602));
   HA_X1 i_603 (.A(n_581), .B(n_596), .CO(n_604), .S(n_603));
   XNOR2_X1 i_604 (.A(n_119), .B(n_96), .ZN(n_605));
   XNOR2_X1 i_605 (.A(n_605), .B(n_73), .ZN(n_606));
   INV_X1 i_606 (.A(n_606), .ZN(n_607));
   OR3_X1 i_607 (.A1(n_609), .A2(n_610), .A3(n_611), .ZN(n_608));
   NOR2_X1 i_608 (.A1(n_96), .A2(n_119), .ZN(n_609));
   NOR2_X1 i_609 (.A1(n_73), .A2(n_119), .ZN(n_610));
   NOR2_X1 i_610 (.A1(n_73), .A2(n_96), .ZN(n_611));
   XNOR2_X1 i_611 (.A(n_50), .B(n_27), .ZN(n_612));
   XNOR2_X1 i_612 (.A(n_612), .B(n_4), .ZN(n_613));
   INV_X1 i_613 (.A(n_613), .ZN(n_614));
   OR3_X1 i_614 (.A1(n_616), .A2(n_617), .A3(n_618), .ZN(n_615));
   NOR2_X1 i_615 (.A1(n_27), .A2(n_50), .ZN(n_616));
   NOR2_X1 i_616 (.A1(n_4), .A2(n_50), .ZN(n_617));
   NOR2_X1 i_617 (.A1(n_4), .A2(n_27), .ZN(n_618));
   FA_X1 i_618 (.A(n_591), .B(n_597), .CI(n_614), .CO(n_620), .S(n_619));
   HA_X1 i_619 (.A(n_607), .B(n_604), .CO(n_622), .S(n_621));
   XNOR2_X1 i_620 (.A(n_143), .B(n_120), .ZN(n_623));
   XNOR2_X1 i_621 (.A(n_623), .B(n_97), .ZN(n_624));
   INV_X1 i_622 (.A(n_624), .ZN(n_625));
   OR3_X1 i_623 (.A1(n_627), .A2(n_628), .A3(n_629), .ZN(n_626));
   NOR2_X1 i_624 (.A1(n_120), .A2(n_143), .ZN(n_627));
   NOR2_X1 i_625 (.A1(n_97), .A2(n_143), .ZN(n_628));
   NOR2_X1 i_626 (.A1(n_97), .A2(n_120), .ZN(n_629));
   XNOR2_X1 i_627 (.A(n_74), .B(n_51), .ZN(n_630));
   XNOR2_X1 i_628 (.A(n_630), .B(n_28), .ZN(n_631));
   INV_X1 i_629 (.A(n_631), .ZN(n_632));
   OR3_X1 i_630 (.A1(n_634), .A2(n_635), .A3(n_636), .ZN(n_633));
   NOR2_X1 i_631 (.A1(n_51), .A2(n_74), .ZN(n_634));
   NOR2_X1 i_632 (.A1(n_28), .A2(n_74), .ZN(n_635));
   NOR2_X1 i_633 (.A1(n_28), .A2(n_51), .ZN(n_636));
   XNOR2_X1 i_634 (.A(n_5), .B(n_615), .ZN(n_637));
   XNOR2_X1 i_635 (.A(n_637), .B(n_608), .ZN(n_638));
   INV_X1 i_636 (.A(n_638), .ZN(n_639));
   NAND3_X1 i_637 (.A1(n_641), .A2(n_643), .A3(n_644), .ZN(n_640));
   NAND2_X1 i_638 (.A1(n_615), .A2(n_642), .ZN(n_641));
   INV_X1 i_639 (.A(n_5), .ZN(n_642));
   NAND2_X1 i_640 (.A1(n_608), .A2(n_642), .ZN(n_643));
   NAND2_X1 i_641 (.A1(n_608), .A2(n_615), .ZN(n_644));
   FA_X1 i_642 (.A(n_632), .B(n_625), .CI(n_639), .CO(n_646), .S(n_645));
   HA_X1 i_643 (.A(n_622), .B(n_620), .CO(n_648), .S(n_647));
   XNOR2_X1 i_644 (.A(n_167), .B(n_144), .ZN(n_649));
   XNOR2_X1 i_645 (.A(n_649), .B(n_121), .ZN(n_650));
   INV_X1 i_646 (.A(n_650), .ZN(n_651));
   OR3_X1 i_647 (.A1(n_653), .A2(n_654), .A3(n_655), .ZN(n_652));
   NOR2_X1 i_648 (.A1(n_144), .A2(n_167), .ZN(n_653));
   NOR2_X1 i_649 (.A1(n_121), .A2(n_167), .ZN(n_654));
   NOR2_X1 i_650 (.A1(n_121), .A2(n_144), .ZN(n_655));
   XNOR2_X1 i_651 (.A(n_98), .B(n_75), .ZN(n_656));
   XNOR2_X1 i_652 (.A(n_656), .B(n_52), .ZN(n_657));
   INV_X1 i_653 (.A(n_657), .ZN(n_658));
   OR3_X1 i_654 (.A1(n_660), .A2(n_661), .A3(n_662), .ZN(n_659));
   NOR2_X1 i_655 (.A1(n_75), .A2(n_98), .ZN(n_660));
   NOR2_X1 i_656 (.A1(n_52), .A2(n_98), .ZN(n_661));
   NOR2_X1 i_657 (.A1(n_52), .A2(n_75), .ZN(n_662));
   XNOR2_X1 i_658 (.A(n_29), .B(n_6), .ZN(n_663));
   XNOR2_X1 i_659 (.A(n_663), .B(n_633), .ZN(n_664));
   NAND3_X1 i_660 (.A1(n_666), .A2(n_667), .A3(n_669), .ZN(n_665));
   OR2_X1 i_661 (.A1(n_6), .A2(n_29), .ZN(n_666));
   NAND2_X1 i_662 (.A1(n_633), .A2(n_668), .ZN(n_667));
   INV_X1 i_663 (.A(n_29), .ZN(n_668));
   NAND2_X1 i_664 (.A1(n_633), .A2(n_670), .ZN(n_669));
   INV_X1 i_665 (.A(n_6), .ZN(n_670));
   FA_X1 i_666 (.A(n_626), .B(n_640), .CI(n_664), .CO(n_672), .S(n_671));
   FA_X1 i_667 (.A(n_658), .B(n_651), .CI(n_648), .CO(n_674), .S(n_673));
   HA_X1 i_668 (.A(n_671), .B(n_646), .CO(n_676), .S(n_675));
   XNOR2_X1 i_669 (.A(n_191), .B(n_168), .ZN(n_677));
   XNOR2_X1 i_670 (.A(n_677), .B(n_145), .ZN(n_678));
   INV_X1 i_671 (.A(n_678), .ZN(n_679));
   OR3_X1 i_672 (.A1(n_681), .A2(n_682), .A3(n_683), .ZN(n_680));
   NOR2_X1 i_673 (.A1(n_168), .A2(n_191), .ZN(n_681));
   NOR2_X1 i_674 (.A1(n_145), .A2(n_191), .ZN(n_682));
   NOR2_X1 i_675 (.A1(n_145), .A2(n_168), .ZN(n_683));
   XNOR2_X1 i_676 (.A(n_122), .B(n_99), .ZN(n_684));
   XNOR2_X1 i_677 (.A(n_684), .B(n_76), .ZN(n_685));
   INV_X1 i_678 (.A(n_685), .ZN(n_686));
   OR3_X1 i_679 (.A1(n_688), .A2(n_689), .A3(n_690), .ZN(n_687));
   NOR2_X1 i_680 (.A1(n_99), .A2(n_122), .ZN(n_688));
   NOR2_X1 i_681 (.A1(n_76), .A2(n_122), .ZN(n_689));
   NOR2_X1 i_682 (.A1(n_76), .A2(n_99), .ZN(n_690));
   XNOR2_X1 i_683 (.A(n_53), .B(n_30), .ZN(n_691));
   XNOR2_X1 i_684 (.A(n_691), .B(n_7), .ZN(n_692));
   INV_X1 i_685 (.A(n_692), .ZN(n_693));
   OR3_X1 i_686 (.A1(n_695), .A2(n_696), .A3(n_697), .ZN(n_694));
   NOR2_X1 i_687 (.A1(n_30), .A2(n_53), .ZN(n_695));
   NOR2_X1 i_688 (.A1(n_7), .A2(n_53), .ZN(n_696));
   NOR2_X1 i_689 (.A1(n_7), .A2(n_30), .ZN(n_697));
   FA_X1 i_690 (.A(n_659), .B(n_652), .CI(n_665), .CO(n_699), .S(n_698));
   FA_X1 i_691 (.A(n_693), .B(n_686), .CI(n_679), .CO(n_701), .S(n_700));
   FA_X1 i_692 (.A(n_698), .B(n_672), .CI(n_676), .CO(n_703), .S(n_702));
   HA_X1 i_693 (.A(n_674), .B(n_700), .CO(n_705), .S(n_704));
   XNOR2_X1 i_694 (.A(n_215), .B(n_192), .ZN(n_706));
   XNOR2_X1 i_695 (.A(n_706), .B(n_169), .ZN(n_707));
   INV_X1 i_696 (.A(n_707), .ZN(n_708));
   OR3_X1 i_697 (.A1(n_710), .A2(n_711), .A3(n_712), .ZN(n_709));
   NOR2_X1 i_698 (.A1(n_192), .A2(n_215), .ZN(n_710));
   NOR2_X1 i_699 (.A1(n_169), .A2(n_215), .ZN(n_711));
   NOR2_X1 i_700 (.A1(n_169), .A2(n_192), .ZN(n_712));
   XNOR2_X1 i_701 (.A(n_146), .B(n_123), .ZN(n_713));
   XNOR2_X1 i_702 (.A(n_713), .B(n_100), .ZN(n_714));
   INV_X1 i_703 (.A(n_714), .ZN(n_715));
   OR3_X1 i_704 (.A1(n_717), .A2(n_718), .A3(n_719), .ZN(n_716));
   NOR2_X1 i_705 (.A1(n_123), .A2(n_146), .ZN(n_717));
   NOR2_X1 i_706 (.A1(n_100), .A2(n_146), .ZN(n_718));
   NOR2_X1 i_707 (.A1(n_100), .A2(n_123), .ZN(n_719));
   XNOR2_X1 i_708 (.A(n_77), .B(n_54), .ZN(n_720));
   XNOR2_X1 i_709 (.A(n_720), .B(n_31), .ZN(n_721));
   INV_X1 i_710 (.A(n_721), .ZN(n_722));
   OR3_X1 i_711 (.A1(n_724), .A2(n_725), .A3(n_726), .ZN(n_723));
   NOR2_X1 i_712 (.A1(n_54), .A2(n_77), .ZN(n_724));
   NOR2_X1 i_713 (.A1(n_31), .A2(n_77), .ZN(n_725));
   NOR2_X1 i_714 (.A1(n_31), .A2(n_54), .ZN(n_726));
   XNOR2_X1 i_715 (.A(n_8), .B(n_694), .ZN(n_727));
   XNOR2_X1 i_716 (.A(n_727), .B(n_687), .ZN(n_728));
   INV_X1 i_717 (.A(n_728), .ZN(n_729));
   NAND3_X1 i_718 (.A1(n_731), .A2(n_733), .A3(n_734), .ZN(n_730));
   NAND2_X1 i_719 (.A1(n_694), .A2(n_732), .ZN(n_731));
   INV_X1 i_720 (.A(n_8), .ZN(n_732));
   NAND2_X1 i_721 (.A1(n_687), .A2(n_732), .ZN(n_733));
   NAND2_X1 i_722 (.A1(n_687), .A2(n_694), .ZN(n_734));
   FA_X1 i_723 (.A(n_680), .B(n_722), .CI(n_715), .CO(n_736), .S(n_735));
   FA_X1 i_724 (.A(n_708), .B(n_699), .CI(n_729), .CO(n_738), .S(n_737));
   FA_X1 i_725 (.A(n_701), .B(n_735), .CI(n_737), .CO(n_740), .S(n_739));
   HA_X1 i_726 (.A(n_705), .B(n_703), .CO(n_742), .S(n_741));
   XNOR2_X1 i_727 (.A(n_239), .B(n_216), .ZN(n_743));
   XNOR2_X1 i_728 (.A(n_743), .B(n_193), .ZN(n_744));
   INV_X1 i_729 (.A(n_744), .ZN(n_745));
   OR3_X1 i_730 (.A1(n_747), .A2(n_748), .A3(n_749), .ZN(n_746));
   NOR2_X1 i_731 (.A1(n_216), .A2(n_239), .ZN(n_747));
   NOR2_X1 i_732 (.A1(n_193), .A2(n_239), .ZN(n_748));
   NOR2_X1 i_733 (.A1(n_193), .A2(n_216), .ZN(n_749));
   XNOR2_X1 i_734 (.A(n_170), .B(n_147), .ZN(n_750));
   XNOR2_X1 i_735 (.A(n_750), .B(n_124), .ZN(n_751));
   INV_X1 i_736 (.A(n_751), .ZN(n_752));
   OR3_X1 i_737 (.A1(n_754), .A2(n_755), .A3(n_756), .ZN(n_753));
   NOR2_X1 i_738 (.A1(n_147), .A2(n_170), .ZN(n_754));
   NOR2_X1 i_739 (.A1(n_124), .A2(n_170), .ZN(n_755));
   NOR2_X1 i_740 (.A1(n_124), .A2(n_147), .ZN(n_756));
   XNOR2_X1 i_741 (.A(n_101), .B(n_78), .ZN(n_757));
   XNOR2_X1 i_742 (.A(n_757), .B(n_55), .ZN(n_758));
   INV_X1 i_743 (.A(n_758), .ZN(n_759));
   OR3_X1 i_744 (.A1(n_761), .A2(n_762), .A3(n_763), .ZN(n_760));
   NOR2_X1 i_745 (.A1(n_78), .A2(n_101), .ZN(n_761));
   NOR2_X1 i_746 (.A1(n_55), .A2(n_101), .ZN(n_762));
   NOR2_X1 i_747 (.A1(n_55), .A2(n_78), .ZN(n_763));
   XNOR2_X1 i_748 (.A(n_32), .B(n_9), .ZN(n_764));
   XNOR2_X1 i_749 (.A(n_764), .B(n_723), .ZN(n_765));
   NAND3_X1 i_750 (.A1(n_767), .A2(n_768), .A3(n_770), .ZN(n_766));
   OR2_X1 i_751 (.A1(n_9), .A2(n_32), .ZN(n_767));
   NAND2_X1 i_752 (.A1(n_723), .A2(n_769), .ZN(n_768));
   INV_X1 i_753 (.A(n_32), .ZN(n_769));
   NAND2_X1 i_754 (.A1(n_723), .A2(n_771), .ZN(n_770));
   INV_X1 i_755 (.A(n_9), .ZN(n_771));
   FA_X1 i_756 (.A(n_716), .B(n_709), .CI(n_730), .CO(n_773), .S(n_772));
   FA_X1 i_757 (.A(n_765), .B(n_759), .CI(n_752), .CO(n_775), .S(n_774));
   FA_X1 i_758 (.A(n_745), .B(n_772), .CI(n_736), .CO(n_777), .S(n_776));
   FA_X1 i_759 (.A(n_738), .B(n_774), .CI(n_776), .CO(n_779), .S(n_778));
   HA_X1 i_760 (.A(n_742), .B(n_740), .CO(n_781), .S(n_780));
   XNOR2_X1 i_761 (.A(n_263), .B(n_240), .ZN(n_782));
   XNOR2_X1 i_762 (.A(n_782), .B(n_217), .ZN(n_783));
   INV_X1 i_763 (.A(n_783), .ZN(n_784));
   OR3_X1 i_764 (.A1(n_786), .A2(n_787), .A3(n_788), .ZN(n_785));
   NOR2_X1 i_765 (.A1(n_240), .A2(n_263), .ZN(n_786));
   NOR2_X1 i_766 (.A1(n_217), .A2(n_263), .ZN(n_787));
   NOR2_X1 i_767 (.A1(n_217), .A2(n_240), .ZN(n_788));
   XNOR2_X1 i_768 (.A(n_194), .B(n_171), .ZN(n_789));
   XNOR2_X1 i_769 (.A(n_789), .B(n_148), .ZN(n_790));
   INV_X1 i_770 (.A(n_790), .ZN(n_791));
   OR3_X1 i_771 (.A1(n_793), .A2(n_794), .A3(n_795), .ZN(n_792));
   NOR2_X1 i_772 (.A1(n_171), .A2(n_194), .ZN(n_793));
   NOR2_X1 i_773 (.A1(n_148), .A2(n_194), .ZN(n_794));
   NOR2_X1 i_774 (.A1(n_148), .A2(n_171), .ZN(n_795));
   XNOR2_X1 i_775 (.A(n_125), .B(n_102), .ZN(n_796));
   XNOR2_X1 i_776 (.A(n_796), .B(n_79), .ZN(n_797));
   INV_X1 i_777 (.A(n_797), .ZN(n_798));
   OR3_X1 i_778 (.A1(n_800), .A2(n_801), .A3(n_802), .ZN(n_799));
   NOR2_X1 i_779 (.A1(n_102), .A2(n_125), .ZN(n_800));
   NOR2_X1 i_780 (.A1(n_79), .A2(n_125), .ZN(n_801));
   NOR2_X1 i_781 (.A1(n_79), .A2(n_102), .ZN(n_802));
   XNOR2_X1 i_782 (.A(n_56), .B(n_33), .ZN(n_803));
   XNOR2_X1 i_783 (.A(n_803), .B(n_10), .ZN(n_804));
   INV_X1 i_784 (.A(n_804), .ZN(n_805));
   OR3_X1 i_785 (.A1(n_807), .A2(n_808), .A3(n_809), .ZN(n_806));
   NOR2_X1 i_786 (.A1(n_33), .A2(n_56), .ZN(n_807));
   NOR2_X1 i_787 (.A1(n_10), .A2(n_56), .ZN(n_808));
   NOR2_X1 i_788 (.A1(n_10), .A2(n_33), .ZN(n_809));
   FA_X1 i_789 (.A(n_760), .B(n_753), .CI(n_746), .CO(n_811), .S(n_810));
   FA_X1 i_790 (.A(n_766), .B(n_805), .CI(n_798), .CO(n_813), .S(n_812));
   FA_X1 i_791 (.A(n_791), .B(n_784), .CI(n_773), .CO(n_815), .S(n_814));
   FA_X1 i_792 (.A(n_810), .B(n_775), .CI(n_777), .CO(n_817), .S(n_816));
   FA_X1 i_793 (.A(n_814), .B(n_812), .CI(n_816), .CO(n_819), .S(n_818));
   HA_X1 i_794 (.A(n_781), .B(n_779), .CO(n_821), .S(n_820));
   XNOR2_X1 i_795 (.A(n_287), .B(n_264), .ZN(n_822));
   XNOR2_X1 i_796 (.A(n_822), .B(n_241), .ZN(n_823));
   INV_X1 i_797 (.A(n_823), .ZN(n_824));
   OR3_X1 i_798 (.A1(n_826), .A2(n_827), .A3(n_828), .ZN(n_825));
   NOR2_X1 i_799 (.A1(n_264), .A2(n_287), .ZN(n_826));
   NOR2_X1 i_800 (.A1(n_241), .A2(n_287), .ZN(n_827));
   NOR2_X1 i_801 (.A1(n_241), .A2(n_264), .ZN(n_828));
   XNOR2_X1 i_802 (.A(n_218), .B(n_195), .ZN(n_829));
   XNOR2_X1 i_803 (.A(n_829), .B(n_172), .ZN(n_830));
   INV_X1 i_804 (.A(n_830), .ZN(n_831));
   OR3_X1 i_805 (.A1(n_833), .A2(n_834), .A3(n_835), .ZN(n_832));
   NOR2_X1 i_806 (.A1(n_195), .A2(n_218), .ZN(n_833));
   NOR2_X1 i_807 (.A1(n_172), .A2(n_218), .ZN(n_834));
   NOR2_X1 i_808 (.A1(n_172), .A2(n_195), .ZN(n_835));
   XNOR2_X1 i_809 (.A(n_149), .B(n_126), .ZN(n_836));
   XNOR2_X1 i_810 (.A(n_836), .B(n_103), .ZN(n_837));
   INV_X1 i_811 (.A(n_837), .ZN(n_838));
   OR3_X1 i_812 (.A1(n_840), .A2(n_841), .A3(n_842), .ZN(n_839));
   NOR2_X1 i_813 (.A1(n_126), .A2(n_149), .ZN(n_840));
   NOR2_X1 i_814 (.A1(n_103), .A2(n_149), .ZN(n_841));
   NOR2_X1 i_815 (.A1(n_103), .A2(n_126), .ZN(n_842));
   XNOR2_X1 i_816 (.A(n_80), .B(n_57), .ZN(n_843));
   XNOR2_X1 i_817 (.A(n_843), .B(n_34), .ZN(n_844));
   INV_X1 i_818 (.A(n_844), .ZN(n_845));
   OR3_X1 i_819 (.A1(n_847), .A2(n_848), .A3(n_849), .ZN(n_846));
   NOR2_X1 i_820 (.A1(n_57), .A2(n_80), .ZN(n_847));
   NOR2_X1 i_821 (.A1(n_34), .A2(n_80), .ZN(n_848));
   NOR2_X1 i_822 (.A1(n_34), .A2(n_57), .ZN(n_849));
   XNOR2_X1 i_823 (.A(n_11), .B(n_806), .ZN(n_850));
   XNOR2_X1 i_824 (.A(n_850), .B(n_799), .ZN(n_851));
   INV_X1 i_825 (.A(n_851), .ZN(n_852));
   NAND3_X1 i_826 (.A1(n_854), .A2(n_856), .A3(n_857), .ZN(n_853));
   NAND2_X1 i_827 (.A1(n_806), .A2(n_855), .ZN(n_854));
   INV_X1 i_828 (.A(n_11), .ZN(n_855));
   NAND2_X1 i_829 (.A1(n_799), .A2(n_855), .ZN(n_856));
   NAND2_X1 i_830 (.A1(n_799), .A2(n_806), .ZN(n_857));
   FA_X1 i_831 (.A(n_792), .B(n_785), .CI(n_811), .CO(n_859), .S(n_858));
   FA_X1 i_832 (.A(n_845), .B(n_838), .CI(n_831), .CO(n_861), .S(n_860));
   FA_X1 i_833 (.A(n_824), .B(n_858), .CI(n_852), .CO(n_863), .S(n_862));
   FA_X1 i_834 (.A(n_813), .B(n_815), .CI(n_860), .CO(n_865), .S(n_864));
   FA_X1 i_835 (.A(n_817), .B(n_862), .CI(n_864), .CO(n_867), .S(n_866));
   HA_X1 i_836 (.A(n_819), .B(n_821), .CO(n_869), .S(n_868));
   XNOR2_X1 i_837 (.A(n_311), .B(n_288), .ZN(n_870));
   XNOR2_X1 i_838 (.A(n_870), .B(n_265), .ZN(n_871));
   INV_X1 i_839 (.A(n_871), .ZN(n_872));
   OR3_X1 i_840 (.A1(n_874), .A2(n_875), .A3(n_876), .ZN(n_873));
   NOR2_X1 i_841 (.A1(n_288), .A2(n_311), .ZN(n_874));
   NOR2_X1 i_842 (.A1(n_265), .A2(n_311), .ZN(n_875));
   NOR2_X1 i_843 (.A1(n_265), .A2(n_288), .ZN(n_876));
   XNOR2_X1 i_844 (.A(n_242), .B(n_219), .ZN(n_877));
   XNOR2_X1 i_845 (.A(n_877), .B(n_196), .ZN(n_878));
   INV_X1 i_846 (.A(n_878), .ZN(n_879));
   OR3_X1 i_847 (.A1(n_881), .A2(n_882), .A3(n_883), .ZN(n_880));
   NOR2_X1 i_848 (.A1(n_219), .A2(n_242), .ZN(n_881));
   NOR2_X1 i_849 (.A1(n_196), .A2(n_242), .ZN(n_882));
   NOR2_X1 i_850 (.A1(n_196), .A2(n_219), .ZN(n_883));
   XNOR2_X1 i_851 (.A(n_173), .B(n_150), .ZN(n_884));
   XNOR2_X1 i_852 (.A(n_884), .B(n_127), .ZN(n_885));
   INV_X1 i_853 (.A(n_885), .ZN(n_886));
   OR3_X1 i_854 (.A1(n_888), .A2(n_889), .A3(n_890), .ZN(n_887));
   NOR2_X1 i_855 (.A1(n_150), .A2(n_173), .ZN(n_888));
   NOR2_X1 i_856 (.A1(n_127), .A2(n_173), .ZN(n_889));
   NOR2_X1 i_857 (.A1(n_127), .A2(n_150), .ZN(n_890));
   XNOR2_X1 i_858 (.A(n_104), .B(n_81), .ZN(n_891));
   XNOR2_X1 i_859 (.A(n_891), .B(n_58), .ZN(n_892));
   INV_X1 i_860 (.A(n_892), .ZN(n_893));
   OR3_X1 i_861 (.A1(n_895), .A2(n_896), .A3(n_897), .ZN(n_894));
   NOR2_X1 i_862 (.A1(n_81), .A2(n_104), .ZN(n_895));
   NOR2_X1 i_863 (.A1(n_58), .A2(n_104), .ZN(n_896));
   NOR2_X1 i_864 (.A1(n_58), .A2(n_81), .ZN(n_897));
   XNOR2_X1 i_865 (.A(n_35), .B(n_12), .ZN(n_898));
   XNOR2_X1 i_866 (.A(n_898), .B(n_846), .ZN(n_899));
   NAND3_X1 i_867 (.A1(n_901), .A2(n_902), .A3(n_904), .ZN(n_900));
   OR2_X1 i_868 (.A1(n_12), .A2(n_35), .ZN(n_901));
   NAND2_X1 i_869 (.A1(n_846), .A2(n_903), .ZN(n_902));
   INV_X1 i_870 (.A(n_35), .ZN(n_903));
   NAND2_X1 i_871 (.A1(n_846), .A2(n_905), .ZN(n_904));
   INV_X1 i_872 (.A(n_12), .ZN(n_905));
   FA_X1 i_873 (.A(n_839), .B(n_832), .CI(n_825), .CO(n_907), .S(n_906));
   FA_X1 i_874 (.A(n_853), .B(n_899), .CI(n_893), .CO(n_909), .S(n_908));
   FA_X1 i_875 (.A(n_886), .B(n_879), .CI(n_872), .CO(n_911), .S(n_910));
   FA_X1 i_876 (.A(n_859), .B(n_906), .CI(n_861), .CO(n_913), .S(n_912));
   FA_X1 i_877 (.A(n_863), .B(n_910), .CI(n_908), .CO(n_915), .S(n_914));
   FA_X1 i_878 (.A(n_912), .B(n_865), .CI(n_867), .CO(n_917), .S(n_916));
   HA_X1 i_879 (.A(n_914), .B(n_869), .CO(n_919), .S(n_918));
   XNOR2_X1 i_880 (.A(n_335), .B(n_312), .ZN(n_920));
   XNOR2_X1 i_881 (.A(n_920), .B(n_289), .ZN(n_921));
   INV_X1 i_882 (.A(n_921), .ZN(n_922));
   OR3_X1 i_883 (.A1(n_924), .A2(n_925), .A3(n_926), .ZN(n_923));
   NOR2_X1 i_884 (.A1(n_312), .A2(n_335), .ZN(n_924));
   NOR2_X1 i_885 (.A1(n_289), .A2(n_335), .ZN(n_925));
   NOR2_X1 i_886 (.A1(n_289), .A2(n_312), .ZN(n_926));
   XNOR2_X1 i_887 (.A(n_266), .B(n_243), .ZN(n_927));
   XNOR2_X1 i_888 (.A(n_927), .B(n_220), .ZN(n_928));
   INV_X1 i_889 (.A(n_928), .ZN(n_929));
   OR3_X1 i_890 (.A1(n_931), .A2(n_932), .A3(n_933), .ZN(n_930));
   NOR2_X1 i_891 (.A1(n_243), .A2(n_266), .ZN(n_931));
   NOR2_X1 i_892 (.A1(n_220), .A2(n_266), .ZN(n_932));
   NOR2_X1 i_893 (.A1(n_220), .A2(n_243), .ZN(n_933));
   XNOR2_X1 i_894 (.A(n_197), .B(n_174), .ZN(n_934));
   XNOR2_X1 i_895 (.A(n_934), .B(n_151), .ZN(n_935));
   INV_X1 i_896 (.A(n_935), .ZN(n_936));
   OR3_X1 i_897 (.A1(n_938), .A2(n_939), .A3(n_940), .ZN(n_937));
   NOR2_X1 i_898 (.A1(n_174), .A2(n_197), .ZN(n_938));
   NOR2_X1 i_899 (.A1(n_151), .A2(n_197), .ZN(n_939));
   NOR2_X1 i_900 (.A1(n_151), .A2(n_174), .ZN(n_940));
   XNOR2_X1 i_901 (.A(n_128), .B(n_105), .ZN(n_941));
   XNOR2_X1 i_902 (.A(n_941), .B(n_82), .ZN(n_942));
   INV_X1 i_903 (.A(n_942), .ZN(n_943));
   OR3_X1 i_904 (.A1(n_945), .A2(n_946), .A3(n_947), .ZN(n_944));
   NOR2_X1 i_905 (.A1(n_105), .A2(n_128), .ZN(n_945));
   NOR2_X1 i_906 (.A1(n_82), .A2(n_128), .ZN(n_946));
   NOR2_X1 i_907 (.A1(n_82), .A2(n_105), .ZN(n_947));
   XNOR2_X1 i_908 (.A(n_59), .B(n_36), .ZN(n_948));
   XNOR2_X1 i_909 (.A(n_948), .B(n_13), .ZN(n_949));
   INV_X1 i_910 (.A(n_949), .ZN(n_950));
   OR3_X1 i_911 (.A1(n_952), .A2(n_953), .A3(n_954), .ZN(n_951));
   NOR2_X1 i_912 (.A1(n_36), .A2(n_59), .ZN(n_952));
   NOR2_X1 i_913 (.A1(n_13), .A2(n_59), .ZN(n_953));
   NOR2_X1 i_914 (.A1(n_13), .A2(n_36), .ZN(n_954));
   FA_X1 i_915 (.A(n_894), .B(n_887), .CI(n_880), .CO(n_956), .S(n_955));
   FA_X1 i_916 (.A(n_873), .B(n_907), .CI(n_900), .CO(n_958), .S(n_957));
   FA_X1 i_917 (.A(n_950), .B(n_943), .CI(n_936), .CO(n_960), .S(n_959));
   FA_X1 i_918 (.A(n_929), .B(n_922), .CI(n_955), .CO(n_962), .S(n_961));
   FA_X1 i_919 (.A(n_911), .B(n_909), .CI(n_957), .CO(n_964), .S(n_963));
   FA_X1 i_920 (.A(n_913), .B(n_961), .CI(n_959), .CO(n_966), .S(n_965));
   FA_X1 i_921 (.A(n_963), .B(n_915), .CI(n_965), .CO(n_968), .S(n_967));
   HA_X1 i_922 (.A(n_917), .B(n_919), .CO(n_970), .S(n_969));
   XNOR2_X1 i_923 (.A(n_359), .B(n_336), .ZN(n_971));
   XNOR2_X1 i_924 (.A(n_971), .B(n_313), .ZN(n_972));
   INV_X1 i_925 (.A(n_972), .ZN(n_973));
   OR3_X1 i_926 (.A1(n_975), .A2(n_976), .A3(n_977), .ZN(n_974));
   NOR2_X1 i_927 (.A1(n_336), .A2(n_359), .ZN(n_975));
   NOR2_X1 i_928 (.A1(n_313), .A2(n_359), .ZN(n_976));
   NOR2_X1 i_929 (.A1(n_313), .A2(n_336), .ZN(n_977));
   XNOR2_X1 i_930 (.A(n_290), .B(n_267), .ZN(n_978));
   XNOR2_X1 i_931 (.A(n_978), .B(n_244), .ZN(n_979));
   INV_X1 i_932 (.A(n_979), .ZN(n_980));
   OR3_X1 i_933 (.A1(n_982), .A2(n_983), .A3(n_984), .ZN(n_981));
   NOR2_X1 i_934 (.A1(n_267), .A2(n_290), .ZN(n_982));
   NOR2_X1 i_935 (.A1(n_244), .A2(n_290), .ZN(n_983));
   NOR2_X1 i_936 (.A1(n_244), .A2(n_267), .ZN(n_984));
   XNOR2_X1 i_937 (.A(n_221), .B(n_198), .ZN(n_985));
   XNOR2_X1 i_938 (.A(n_985), .B(n_175), .ZN(n_986));
   INV_X1 i_939 (.A(n_986), .ZN(n_987));
   OR3_X1 i_940 (.A1(n_989), .A2(n_990), .A3(n_991), .ZN(n_988));
   NOR2_X1 i_941 (.A1(n_198), .A2(n_221), .ZN(n_989));
   NOR2_X1 i_942 (.A1(n_175), .A2(n_221), .ZN(n_990));
   NOR2_X1 i_943 (.A1(n_175), .A2(n_198), .ZN(n_991));
   XNOR2_X1 i_944 (.A(n_152), .B(n_129), .ZN(n_992));
   XNOR2_X1 i_945 (.A(n_992), .B(n_106), .ZN(n_993));
   INV_X1 i_946 (.A(n_993), .ZN(n_994));
   OR3_X1 i_947 (.A1(n_996), .A2(n_997), .A3(n_998), .ZN(n_995));
   NOR2_X1 i_948 (.A1(n_129), .A2(n_152), .ZN(n_996));
   NOR2_X1 i_949 (.A1(n_106), .A2(n_152), .ZN(n_997));
   NOR2_X1 i_950 (.A1(n_106), .A2(n_129), .ZN(n_998));
   XNOR2_X1 i_951 (.A(n_83), .B(n_60), .ZN(n_999));
   XNOR2_X1 i_952 (.A(n_999), .B(n_37), .ZN(n_1000));
   INV_X1 i_953 (.A(n_1000), .ZN(n_1001));
   OR3_X1 i_954 (.A1(n_1003), .A2(n_1004), .A3(n_1005), .ZN(n_1002));
   NOR2_X1 i_955 (.A1(n_60), .A2(n_83), .ZN(n_1003));
   NOR2_X1 i_956 (.A1(n_37), .A2(n_83), .ZN(n_1004));
   NOR2_X1 i_957 (.A1(n_37), .A2(n_60), .ZN(n_1005));
   XNOR2_X1 i_958 (.A(n_14), .B(n_951), .ZN(n_1006));
   XNOR2_X1 i_959 (.A(n_1006), .B(n_944), .ZN(n_1007));
   INV_X1 i_960 (.A(n_1007), .ZN(n_1008));
   NAND3_X1 i_961 (.A1(n_1010), .A2(n_1012), .A3(n_1013), .ZN(n_1009));
   NAND2_X1 i_962 (.A1(n_951), .A2(n_1011), .ZN(n_1010));
   INV_X1 i_963 (.A(n_14), .ZN(n_1011));
   NAND2_X1 i_964 (.A1(n_944), .A2(n_1011), .ZN(n_1012));
   NAND2_X1 i_965 (.A1(n_944), .A2(n_951), .ZN(n_1013));
   FA_X1 i_966 (.A(n_937), .B(n_930), .CI(n_923), .CO(n_1015), .S(n_1014));
   FA_X1 i_967 (.A(n_956), .B(n_1001), .CI(n_994), .CO(n_1017), .S(n_1016));
   FA_X1 i_968 (.A(n_987), .B(n_980), .CI(n_973), .CO(n_1019), .S(n_1018));
   FA_X1 i_969 (.A(n_958), .B(n_1014), .CI(n_1008), .CO(n_1021), .S(n_1020));
   FA_X1 i_970 (.A(n_960), .B(n_962), .CI(n_1018), .CO(n_1023), .S(n_1022));
   FA_X1 i_971 (.A(n_1016), .B(n_964), .CI(n_1020), .CO(n_1025), .S(n_1024));
   FA_X1 i_972 (.A(n_966), .B(n_1022), .CI(n_1024), .CO(n_1027), .S(n_1026));
   HA_X1 i_973 (.A(n_968), .B(n_970), .CO(n_1029), .S(n_1028));
   XNOR2_X1 i_974 (.A(n_383), .B(n_360), .ZN(n_1030));
   XNOR2_X1 i_975 (.A(n_1030), .B(n_337), .ZN(n_1031));
   INV_X1 i_976 (.A(n_1031), .ZN(n_1032));
   OR3_X1 i_977 (.A1(n_1034), .A2(n_1035), .A3(n_1036), .ZN(n_1033));
   NOR2_X1 i_978 (.A1(n_360), .A2(n_383), .ZN(n_1034));
   NOR2_X1 i_979 (.A1(n_337), .A2(n_383), .ZN(n_1035));
   NOR2_X1 i_980 (.A1(n_337), .A2(n_360), .ZN(n_1036));
   XNOR2_X1 i_981 (.A(n_314), .B(n_291), .ZN(n_1037));
   XNOR2_X1 i_982 (.A(n_1037), .B(n_268), .ZN(n_1038));
   INV_X1 i_983 (.A(n_1038), .ZN(n_1039));
   OR3_X1 i_984 (.A1(n_1041), .A2(n_1042), .A3(n_1043), .ZN(n_1040));
   NOR2_X1 i_985 (.A1(n_291), .A2(n_314), .ZN(n_1041));
   NOR2_X1 i_986 (.A1(n_268), .A2(n_314), .ZN(n_1042));
   NOR2_X1 i_987 (.A1(n_268), .A2(n_291), .ZN(n_1043));
   XNOR2_X1 i_988 (.A(n_245), .B(n_222), .ZN(n_1044));
   XNOR2_X1 i_989 (.A(n_1044), .B(n_199), .ZN(n_1045));
   INV_X1 i_990 (.A(n_1045), .ZN(n_1046));
   OR3_X1 i_991 (.A1(n_1048), .A2(n_1049), .A3(n_1050), .ZN(n_1047));
   NOR2_X1 i_992 (.A1(n_222), .A2(n_245), .ZN(n_1048));
   NOR2_X1 i_993 (.A1(n_199), .A2(n_245), .ZN(n_1049));
   NOR2_X1 i_994 (.A1(n_199), .A2(n_222), .ZN(n_1050));
   XNOR2_X1 i_995 (.A(n_176), .B(n_153), .ZN(n_1051));
   XNOR2_X1 i_996 (.A(n_1051), .B(n_130), .ZN(n_1052));
   INV_X1 i_997 (.A(n_1052), .ZN(n_1053));
   OR3_X1 i_998 (.A1(n_1055), .A2(n_1056), .A3(n_1057), .ZN(n_1054));
   NOR2_X1 i_999 (.A1(n_153), .A2(n_176), .ZN(n_1055));
   NOR2_X1 i_1000 (.A1(n_130), .A2(n_176), .ZN(n_1056));
   NOR2_X1 i_1001 (.A1(n_130), .A2(n_153), .ZN(n_1057));
   XNOR2_X1 i_1002 (.A(n_107), .B(n_84), .ZN(n_1058));
   XNOR2_X1 i_1003 (.A(n_1058), .B(n_61), .ZN(n_1059));
   INV_X1 i_1004 (.A(n_1059), .ZN(n_1060));
   OR3_X1 i_1005 (.A1(n_1062), .A2(n_1063), .A3(n_1064), .ZN(n_1061));
   NOR2_X1 i_1006 (.A1(n_84), .A2(n_107), .ZN(n_1062));
   NOR2_X1 i_1007 (.A1(n_61), .A2(n_107), .ZN(n_1063));
   NOR2_X1 i_1008 (.A1(n_61), .A2(n_84), .ZN(n_1064));
   XNOR2_X1 i_1009 (.A(n_38), .B(n_15), .ZN(n_1065));
   XNOR2_X1 i_1010 (.A(n_1065), .B(n_1002), .ZN(n_1066));
   NAND3_X1 i_1011 (.A1(n_1068), .A2(n_1069), .A3(n_1071), .ZN(n_1067));
   OR2_X1 i_1012 (.A1(n_15), .A2(n_38), .ZN(n_1068));
   NAND2_X1 i_1013 (.A1(n_1002), .A2(n_1070), .ZN(n_1069));
   INV_X1 i_1014 (.A(n_38), .ZN(n_1070));
   NAND2_X1 i_1015 (.A1(n_1002), .A2(n_1072), .ZN(n_1071));
   INV_X1 i_1016 (.A(n_15), .ZN(n_1072));
   FA_X1 i_1017 (.A(n_995), .B(n_988), .CI(n_981), .CO(n_1074), .S(n_1073));
   FA_X1 i_1018 (.A(n_974), .B(n_1015), .CI(n_1009), .CO(n_1076), .S(n_1075));
   FA_X1 i_1019 (.A(n_1066), .B(n_1060), .CI(n_1053), .CO(n_1078), .S(n_1077));
   FA_X1 i_1020 (.A(n_1046), .B(n_1039), .CI(n_1032), .CO(n_1080), .S(n_1079));
   FA_X1 i_1021 (.A(n_1073), .B(n_1019), .CI(n_1017), .CO(n_1082), .S(n_1081));
   FA_X1 i_1022 (.A(n_1075), .B(n_1021), .CI(n_1079), .CO(n_1084), .S(n_1083));
   FA_X1 i_1023 (.A(n_1077), .B(n_1081), .CI(n_1023), .CO(n_1086), .S(n_1085));
   FA_X1 i_1024 (.A(n_1083), .B(n_1025), .CI(n_1085), .CO(n_1088), .S(n_1087));
   HA_X1 i_1025 (.A(n_1027), .B(n_1029), .CO(n_1090), .S(n_1089));
   XNOR2_X1 i_1026 (.A(n_407), .B(n_384), .ZN(n_1091));
   XNOR2_X1 i_1027 (.A(n_1091), .B(n_361), .ZN(n_1092));
   INV_X1 i_1028 (.A(n_1092), .ZN(n_1093));
   OR3_X1 i_1029 (.A1(n_1095), .A2(n_1096), .A3(n_1097), .ZN(n_1094));
   NOR2_X1 i_1030 (.A1(n_384), .A2(n_407), .ZN(n_1095));
   NOR2_X1 i_1031 (.A1(n_361), .A2(n_407), .ZN(n_1096));
   NOR2_X1 i_1032 (.A1(n_361), .A2(n_384), .ZN(n_1097));
   XNOR2_X1 i_1033 (.A(n_338), .B(n_315), .ZN(n_1098));
   XNOR2_X1 i_1034 (.A(n_1098), .B(n_292), .ZN(n_1099));
   INV_X1 i_1035 (.A(n_1099), .ZN(n_1100));
   OR3_X1 i_1036 (.A1(n_1102), .A2(n_1103), .A3(n_1104), .ZN(n_1101));
   NOR2_X1 i_1037 (.A1(n_315), .A2(n_338), .ZN(n_1102));
   NOR2_X1 i_1038 (.A1(n_292), .A2(n_338), .ZN(n_1103));
   NOR2_X1 i_1039 (.A1(n_292), .A2(n_315), .ZN(n_1104));
   XNOR2_X1 i_1040 (.A(n_269), .B(n_246), .ZN(n_1105));
   XNOR2_X1 i_1041 (.A(n_1105), .B(n_223), .ZN(n_1106));
   INV_X1 i_1042 (.A(n_1106), .ZN(n_1107));
   OR3_X1 i_1043 (.A1(n_1109), .A2(n_1110), .A3(n_1111), .ZN(n_1108));
   NOR2_X1 i_1044 (.A1(n_246), .A2(n_269), .ZN(n_1109));
   NOR2_X1 i_1045 (.A1(n_223), .A2(n_269), .ZN(n_1110));
   NOR2_X1 i_1046 (.A1(n_223), .A2(n_246), .ZN(n_1111));
   XNOR2_X1 i_1047 (.A(n_200), .B(n_177), .ZN(n_1112));
   XNOR2_X1 i_1048 (.A(n_1112), .B(n_154), .ZN(n_1113));
   INV_X1 i_1049 (.A(n_1113), .ZN(n_1114));
   OR3_X1 i_1050 (.A1(n_1116), .A2(n_1117), .A3(n_1118), .ZN(n_1115));
   NOR2_X1 i_1051 (.A1(n_177), .A2(n_200), .ZN(n_1116));
   NOR2_X1 i_1052 (.A1(n_154), .A2(n_200), .ZN(n_1117));
   NOR2_X1 i_1053 (.A1(n_154), .A2(n_177), .ZN(n_1118));
   XNOR2_X1 i_1054 (.A(n_131), .B(n_108), .ZN(n_1119));
   XNOR2_X1 i_1055 (.A(n_1119), .B(n_85), .ZN(n_1120));
   INV_X1 i_1056 (.A(n_1120), .ZN(n_1121));
   OR3_X1 i_1057 (.A1(n_1123), .A2(n_1124), .A3(n_1125), .ZN(n_1122));
   NOR2_X1 i_1058 (.A1(n_108), .A2(n_131), .ZN(n_1123));
   NOR2_X1 i_1059 (.A1(n_85), .A2(n_131), .ZN(n_1124));
   NOR2_X1 i_1060 (.A1(n_85), .A2(n_108), .ZN(n_1125));
   XNOR2_X1 i_1061 (.A(n_62), .B(n_39), .ZN(n_1126));
   XNOR2_X1 i_1062 (.A(n_1126), .B(n_16), .ZN(n_1127));
   INV_X1 i_1063 (.A(n_1127), .ZN(n_1128));
   OR3_X1 i_1064 (.A1(n_1130), .A2(n_1131), .A3(n_1132), .ZN(n_1129));
   NOR2_X1 i_1065 (.A1(n_39), .A2(n_62), .ZN(n_1130));
   NOR2_X1 i_1066 (.A1(n_16), .A2(n_62), .ZN(n_1131));
   NOR2_X1 i_1067 (.A1(n_16), .A2(n_39), .ZN(n_1132));
   FA_X1 i_1068 (.A(n_1061), .B(n_1054), .CI(n_1047), .CO(n_1134), .S(n_1133));
   FA_X1 i_1069 (.A(n_1040), .B(n_1033), .CI(n_1074), .CO(n_1136), .S(n_1135));
   FA_X1 i_1070 (.A(n_1067), .B(n_1128), .CI(n_1121), .CO(n_1138), .S(n_1137));
   FA_X1 i_1071 (.A(n_1114), .B(n_1107), .CI(n_1100), .CO(n_1140), .S(n_1139));
   FA_X1 i_1072 (.A(n_1093), .B(n_1076), .CI(n_1135), .CO(n_1142), .S(n_1141));
   FA_X1 i_1073 (.A(n_1133), .B(n_1080), .CI(n_1078), .CO(n_1144), .S(n_1143));
   FA_X1 i_1074 (.A(n_1082), .B(n_1139), .CI(n_1137), .CO(n_1146), .S(n_1145));
   FA_X1 i_1075 (.A(n_1141), .B(n_1143), .CI(n_1084), .CO(n_1148), .S(n_1147));
   FA_X1 i_1076 (.A(n_1086), .B(n_1145), .CI(n_1147), .CO(n_1150), .S(n_1149));
   HA_X1 i_1077 (.A(n_1088), .B(n_1090), .CO(n_1152), .S(n_1151));
   XNOR2_X1 i_1078 (.A(n_431), .B(n_408), .ZN(n_1153));
   XNOR2_X1 i_1079 (.A(n_1153), .B(n_385), .ZN(n_1154));
   INV_X1 i_1080 (.A(n_1154), .ZN(n_1155));
   OR3_X1 i_1081 (.A1(n_1157), .A2(n_1158), .A3(n_1159), .ZN(n_1156));
   NOR2_X1 i_1082 (.A1(n_408), .A2(n_431), .ZN(n_1157));
   NOR2_X1 i_1083 (.A1(n_385), .A2(n_431), .ZN(n_1158));
   NOR2_X1 i_1084 (.A1(n_385), .A2(n_408), .ZN(n_1159));
   XNOR2_X1 i_1085 (.A(n_362), .B(n_339), .ZN(n_1160));
   XNOR2_X1 i_1086 (.A(n_1160), .B(n_316), .ZN(n_1161));
   INV_X1 i_1087 (.A(n_1161), .ZN(n_1162));
   OR3_X1 i_1088 (.A1(n_1164), .A2(n_1165), .A3(n_1166), .ZN(n_1163));
   NOR2_X1 i_1089 (.A1(n_339), .A2(n_362), .ZN(n_1164));
   NOR2_X1 i_1090 (.A1(n_316), .A2(n_362), .ZN(n_1165));
   NOR2_X1 i_1091 (.A1(n_316), .A2(n_339), .ZN(n_1166));
   XNOR2_X1 i_1092 (.A(n_293), .B(n_270), .ZN(n_1167));
   XNOR2_X1 i_1093 (.A(n_1167), .B(n_247), .ZN(n_1168));
   INV_X1 i_1094 (.A(n_1168), .ZN(n_1169));
   OR3_X1 i_1095 (.A1(n_1171), .A2(n_1172), .A3(n_1173), .ZN(n_1170));
   NOR2_X1 i_1096 (.A1(n_270), .A2(n_293), .ZN(n_1171));
   NOR2_X1 i_1097 (.A1(n_247), .A2(n_293), .ZN(n_1172));
   NOR2_X1 i_1098 (.A1(n_247), .A2(n_270), .ZN(n_1173));
   XNOR2_X1 i_1099 (.A(n_224), .B(n_201), .ZN(n_1174));
   XNOR2_X1 i_1100 (.A(n_1174), .B(n_178), .ZN(n_1175));
   INV_X1 i_1101 (.A(n_1175), .ZN(n_1176));
   OR3_X1 i_1102 (.A1(n_1178), .A2(n_1179), .A3(n_1180), .ZN(n_1177));
   NOR2_X1 i_1103 (.A1(n_201), .A2(n_224), .ZN(n_1178));
   NOR2_X1 i_1104 (.A1(n_178), .A2(n_224), .ZN(n_1179));
   NOR2_X1 i_1105 (.A1(n_178), .A2(n_201), .ZN(n_1180));
   XNOR2_X1 i_1106 (.A(n_155), .B(n_132), .ZN(n_1181));
   XNOR2_X1 i_1107 (.A(n_1181), .B(n_109), .ZN(n_1182));
   INV_X1 i_1108 (.A(n_1182), .ZN(n_1183));
   OR3_X1 i_1109 (.A1(n_1185), .A2(n_1186), .A3(n_1187), .ZN(n_1184));
   NOR2_X1 i_1110 (.A1(n_132), .A2(n_155), .ZN(n_1185));
   NOR2_X1 i_1111 (.A1(n_109), .A2(n_155), .ZN(n_1186));
   NOR2_X1 i_1112 (.A1(n_109), .A2(n_132), .ZN(n_1187));
   XNOR2_X1 i_1113 (.A(n_86), .B(n_63), .ZN(n_1188));
   XNOR2_X1 i_1114 (.A(n_1188), .B(n_40), .ZN(n_1189));
   INV_X1 i_1115 (.A(n_1189), .ZN(n_1190));
   OR3_X1 i_1116 (.A1(n_1192), .A2(n_1193), .A3(n_1194), .ZN(n_1191));
   NOR2_X1 i_1117 (.A1(n_63), .A2(n_86), .ZN(n_1192));
   NOR2_X1 i_1118 (.A1(n_40), .A2(n_86), .ZN(n_1193));
   NOR2_X1 i_1119 (.A1(n_40), .A2(n_63), .ZN(n_1194));
   XNOR2_X1 i_1120 (.A(n_17), .B(n_1129), .ZN(n_1195));
   XNOR2_X1 i_1121 (.A(n_1195), .B(n_1122), .ZN(n_1196));
   INV_X1 i_1122 (.A(n_1196), .ZN(n_1197));
   NAND3_X1 i_1123 (.A1(n_1199), .A2(n_1201), .A3(n_1202), .ZN(n_1198));
   NAND2_X1 i_1124 (.A1(n_1129), .A2(n_1200), .ZN(n_1199));
   INV_X1 i_1125 (.A(n_17), .ZN(n_1200));
   NAND2_X1 i_1126 (.A1(n_1122), .A2(n_1200), .ZN(n_1201));
   NAND2_X1 i_1127 (.A1(n_1122), .A2(n_1129), .ZN(n_1202));
   FA_X1 i_1128 (.A(n_1115), .B(n_1108), .CI(n_1101), .CO(n_1204), .S(n_1203));
   FA_X1 i_1129 (.A(n_1094), .B(n_1134), .CI(n_1190), .CO(n_1206), .S(n_1205));
   FA_X1 i_1130 (.A(n_1183), .B(n_1176), .CI(n_1169), .CO(n_1208), .S(n_1207));
   FA_X1 i_1131 (.A(n_1162), .B(n_1155), .CI(n_1136), .CO(n_1210), .S(n_1209));
   FA_X1 i_1132 (.A(n_1203), .B(n_1197), .CI(n_1140), .CO(n_1212), .S(n_1211));
   FA_X1 i_1133 (.A(n_1138), .B(n_1205), .CI(n_1144), .CO(n_1214), .S(n_1213));
   FA_X1 i_1134 (.A(n_1142), .B(n_1209), .CI(n_1207), .CO(n_1216), .S(n_1215));
   FA_X1 i_1135 (.A(n_1211), .B(n_1146), .CI(n_1213), .CO(n_1218), .S(n_1217));
   FA_X1 i_1136 (.A(n_1148), .B(n_1215), .CI(n_1217), .CO(n_1220), .S(n_1219));
   HA_X1 i_1137 (.A(n_1150), .B(n_1219), .CO(n_1222), .S(n_1221));
   XNOR2_X1 i_1138 (.A(n_455), .B(n_432), .ZN(n_1223));
   XNOR2_X1 i_1139 (.A(n_1223), .B(n_409), .ZN(n_1224));
   INV_X1 i_1140 (.A(n_1224), .ZN(n_1225));
   OR3_X1 i_1141 (.A1(n_1227), .A2(n_1228), .A3(n_1229), .ZN(n_1226));
   NOR2_X1 i_1142 (.A1(n_432), .A2(n_455), .ZN(n_1227));
   NOR2_X1 i_1143 (.A1(n_409), .A2(n_455), .ZN(n_1228));
   NOR2_X1 i_1144 (.A1(n_409), .A2(n_432), .ZN(n_1229));
   XNOR2_X1 i_1145 (.A(n_386), .B(n_363), .ZN(n_1230));
   XNOR2_X1 i_1146 (.A(n_1230), .B(n_340), .ZN(n_1231));
   INV_X1 i_1147 (.A(n_1231), .ZN(n_1232));
   OR3_X1 i_1148 (.A1(n_1234), .A2(n_1235), .A3(n_1236), .ZN(n_1233));
   NOR2_X1 i_1149 (.A1(n_363), .A2(n_386), .ZN(n_1234));
   NOR2_X1 i_1150 (.A1(n_340), .A2(n_386), .ZN(n_1235));
   NOR2_X1 i_1151 (.A1(n_340), .A2(n_363), .ZN(n_1236));
   XNOR2_X1 i_1152 (.A(n_317), .B(n_294), .ZN(n_1237));
   XNOR2_X1 i_1153 (.A(n_1237), .B(n_271), .ZN(n_1238));
   INV_X1 i_1154 (.A(n_1238), .ZN(n_1239));
   OR3_X1 i_1155 (.A1(n_1241), .A2(n_1242), .A3(n_1243), .ZN(n_1240));
   NOR2_X1 i_1156 (.A1(n_294), .A2(n_317), .ZN(n_1241));
   NOR2_X1 i_1157 (.A1(n_271), .A2(n_317), .ZN(n_1242));
   NOR2_X1 i_1158 (.A1(n_271), .A2(n_294), .ZN(n_1243));
   XNOR2_X1 i_1159 (.A(n_248), .B(n_225), .ZN(n_1244));
   XNOR2_X1 i_1160 (.A(n_1244), .B(n_202), .ZN(n_1245));
   INV_X1 i_1161 (.A(n_1245), .ZN(n_1246));
   OR3_X1 i_1162 (.A1(n_1248), .A2(n_1249), .A3(n_1250), .ZN(n_1247));
   NOR2_X1 i_1163 (.A1(n_225), .A2(n_248), .ZN(n_1248));
   NOR2_X1 i_1164 (.A1(n_202), .A2(n_248), .ZN(n_1249));
   NOR2_X1 i_1165 (.A1(n_202), .A2(n_225), .ZN(n_1250));
   XNOR2_X1 i_1166 (.A(n_179), .B(n_156), .ZN(n_1251));
   XNOR2_X1 i_1167 (.A(n_1251), .B(n_133), .ZN(n_1252));
   INV_X1 i_1168 (.A(n_1252), .ZN(n_1253));
   OR3_X1 i_1169 (.A1(n_1255), .A2(n_1256), .A3(n_1257), .ZN(n_1254));
   NOR2_X1 i_1170 (.A1(n_156), .A2(n_179), .ZN(n_1255));
   NOR2_X1 i_1171 (.A1(n_133), .A2(n_179), .ZN(n_1256));
   NOR2_X1 i_1172 (.A1(n_133), .A2(n_156), .ZN(n_1257));
   XNOR2_X1 i_1173 (.A(n_110), .B(n_87), .ZN(n_1258));
   XNOR2_X1 i_1174 (.A(n_1258), .B(n_64), .ZN(n_1259));
   INV_X1 i_1175 (.A(n_1259), .ZN(n_1260));
   OR3_X1 i_1176 (.A1(n_1262), .A2(n_1263), .A3(n_1264), .ZN(n_1261));
   NOR2_X1 i_1177 (.A1(n_87), .A2(n_110), .ZN(n_1262));
   NOR2_X1 i_1178 (.A1(n_64), .A2(n_110), .ZN(n_1263));
   NOR2_X1 i_1179 (.A1(n_64), .A2(n_87), .ZN(n_1264));
   XNOR2_X1 i_1180 (.A(n_41), .B(n_18), .ZN(n_1265));
   XNOR2_X1 i_1181 (.A(n_1265), .B(n_1191), .ZN(n_1266));
   NAND3_X1 i_1182 (.A1(n_1268), .A2(n_1269), .A3(n_1271), .ZN(n_1267));
   OR2_X1 i_1183 (.A1(n_18), .A2(n_41), .ZN(n_1268));
   NAND2_X1 i_1184 (.A1(n_1191), .A2(n_1270), .ZN(n_1269));
   INV_X1 i_1185 (.A(n_41), .ZN(n_1270));
   NAND2_X1 i_1186 (.A1(n_1191), .A2(n_1272), .ZN(n_1271));
   INV_X1 i_1187 (.A(n_18), .ZN(n_1272));
   FA_X1 i_1188 (.A(n_1184), .B(n_1177), .CI(n_1170), .CO(n_1274), .S(n_1273));
   FA_X1 i_1189 (.A(n_1163), .B(n_1156), .CI(n_1204), .CO(n_1276), .S(n_1275));
   FA_X1 i_1190 (.A(n_1198), .B(n_1266), .CI(n_1260), .CO(n_1278), .S(n_1277));
   FA_X1 i_1191 (.A(n_1253), .B(n_1246), .CI(n_1239), .CO(n_1280), .S(n_1279));
   FA_X1 i_1192 (.A(n_1232), .B(n_1225), .CI(n_1275), .CO(n_1282), .S(n_1281));
   FA_X1 i_1193 (.A(n_1273), .B(n_1208), .CI(n_1206), .CO(n_1284), .S(n_1283));
   FA_X1 i_1194 (.A(n_1210), .B(n_1212), .CI(n_1281), .CO(n_1286), .S(n_1285));
   FA_X1 i_1195 (.A(n_1279), .B(n_1277), .CI(n_1214), .CO(n_1288), .S(n_1287));
   FA_X1 i_1196 (.A(n_1283), .B(n_1216), .CI(n_1285), .CO(n_1290), .S(n_1289));
   FA_X1 i_1197 (.A(n_1287), .B(n_1218), .CI(n_1289), .CO(n_1292), .S(n_1291));
   HA_X1 i_1198 (.A(n_1220), .B(n_1291), .CO(n_1294), .S(n_1293));
   XNOR2_X1 i_1199 (.A(n_479), .B(n_456), .ZN(n_1295));
   XNOR2_X1 i_1200 (.A(n_1295), .B(n_433), .ZN(n_1296));
   INV_X1 i_1201 (.A(n_1296), .ZN(n_1297));
   OR3_X1 i_1202 (.A1(n_1299), .A2(n_1300), .A3(n_1301), .ZN(n_1298));
   NOR2_X1 i_1203 (.A1(n_456), .A2(n_479), .ZN(n_1299));
   NOR2_X1 i_1204 (.A1(n_433), .A2(n_479), .ZN(n_1300));
   NOR2_X1 i_1205 (.A1(n_433), .A2(n_456), .ZN(n_1301));
   XNOR2_X1 i_1206 (.A(n_410), .B(n_387), .ZN(n_1302));
   XNOR2_X1 i_1207 (.A(n_1302), .B(n_364), .ZN(n_1303));
   INV_X1 i_1208 (.A(n_1303), .ZN(n_1304));
   OR3_X1 i_1209 (.A1(n_1306), .A2(n_1307), .A3(n_1308), .ZN(n_1305));
   NOR2_X1 i_1210 (.A1(n_387), .A2(n_410), .ZN(n_1306));
   NOR2_X1 i_1211 (.A1(n_364), .A2(n_410), .ZN(n_1307));
   NOR2_X1 i_1212 (.A1(n_364), .A2(n_387), .ZN(n_1308));
   XNOR2_X1 i_1213 (.A(n_341), .B(n_318), .ZN(n_1309));
   XNOR2_X1 i_1214 (.A(n_1309), .B(n_295), .ZN(n_1310));
   INV_X1 i_1215 (.A(n_1310), .ZN(n_1311));
   OR3_X1 i_1216 (.A1(n_1313), .A2(n_1314), .A3(n_1315), .ZN(n_1312));
   NOR2_X1 i_1217 (.A1(n_318), .A2(n_341), .ZN(n_1313));
   NOR2_X1 i_1218 (.A1(n_295), .A2(n_341), .ZN(n_1314));
   NOR2_X1 i_1219 (.A1(n_295), .A2(n_318), .ZN(n_1315));
   XNOR2_X1 i_1220 (.A(n_272), .B(n_249), .ZN(n_1316));
   XNOR2_X1 i_1221 (.A(n_1316), .B(n_226), .ZN(n_1317));
   INV_X1 i_1222 (.A(n_1317), .ZN(n_1318));
   OR3_X1 i_1223 (.A1(n_1320), .A2(n_1321), .A3(n_1322), .ZN(n_1319));
   NOR2_X1 i_1224 (.A1(n_249), .A2(n_272), .ZN(n_1320));
   NOR2_X1 i_1225 (.A1(n_226), .A2(n_272), .ZN(n_1321));
   NOR2_X1 i_1226 (.A1(n_226), .A2(n_249), .ZN(n_1322));
   XNOR2_X1 i_1227 (.A(n_203), .B(n_180), .ZN(n_1323));
   XNOR2_X1 i_1228 (.A(n_1323), .B(n_157), .ZN(n_1324));
   INV_X1 i_1229 (.A(n_1324), .ZN(n_1325));
   OR3_X1 i_1230 (.A1(n_1327), .A2(n_1328), .A3(n_1329), .ZN(n_1326));
   NOR2_X1 i_1231 (.A1(n_180), .A2(n_203), .ZN(n_1327));
   NOR2_X1 i_1232 (.A1(n_157), .A2(n_203), .ZN(n_1328));
   NOR2_X1 i_1233 (.A1(n_157), .A2(n_180), .ZN(n_1329));
   XNOR2_X1 i_1234 (.A(n_134), .B(n_111), .ZN(n_1330));
   XNOR2_X1 i_1235 (.A(n_1330), .B(n_88), .ZN(n_1331));
   INV_X1 i_1236 (.A(n_1331), .ZN(n_1332));
   OR3_X1 i_1237 (.A1(n_1334), .A2(n_1335), .A3(n_1336), .ZN(n_1333));
   NOR2_X1 i_1238 (.A1(n_111), .A2(n_134), .ZN(n_1334));
   NOR2_X1 i_1239 (.A1(n_88), .A2(n_134), .ZN(n_1335));
   NOR2_X1 i_1240 (.A1(n_88), .A2(n_111), .ZN(n_1336));
   XNOR2_X1 i_1241 (.A(n_65), .B(n_42), .ZN(n_1337));
   XNOR2_X1 i_1242 (.A(n_1337), .B(n_19), .ZN(n_1338));
   INV_X1 i_1243 (.A(n_1338), .ZN(n_1339));
   OR3_X1 i_1244 (.A1(n_1341), .A2(n_1342), .A3(n_1343), .ZN(n_1340));
   NOR2_X1 i_1245 (.A1(n_42), .A2(n_65), .ZN(n_1341));
   NOR2_X1 i_1246 (.A1(n_19), .A2(n_65), .ZN(n_1342));
   NOR2_X1 i_1247 (.A1(n_19), .A2(n_42), .ZN(n_1343));
   FA_X1 i_1248 (.A(n_1261), .B(n_1254), .CI(n_1247), .CO(n_1345), .S(n_1344));
   FA_X1 i_1249 (.A(n_1240), .B(n_1233), .CI(n_1226), .CO(n_1347), .S(n_1346));
   FA_X1 i_1250 (.A(n_1274), .B(n_1267), .CI(n_1339), .CO(n_1349), .S(n_1348));
   FA_X1 i_1251 (.A(n_1332), .B(n_1325), .CI(n_1318), .CO(n_1351), .S(n_1350));
   FA_X1 i_1252 (.A(n_1311), .B(n_1304), .CI(n_1297), .CO(n_1353), .S(n_1352));
   FA_X1 i_1253 (.A(n_1276), .B(n_1346), .CI(n_1344), .CO(n_1355), .S(n_1354));
   FA_X1 i_1254 (.A(n_1280), .B(n_1278), .CI(n_1348), .CO(n_1357), .S(n_1356));
   FA_X1 i_1255 (.A(n_1284), .B(n_1282), .CI(n_1352), .CO(n_1359), .S(n_1358));
   FA_X1 i_1256 (.A(n_1350), .B(n_1356), .CI(n_1354), .CO(n_1361), .S(n_1360));
   FA_X1 i_1257 (.A(n_1286), .B(n_1288), .CI(n_1358), .CO(n_1363), .S(n_1362));
   FA_X1 i_1258 (.A(n_1290), .B(n_1360), .CI(n_1362), .CO(n_1365), .S(n_1364));
   HA_X1 i_1259 (.A(n_1292), .B(n_1294), .CO(n_1367), .S(n_1366));
   XNOR2_X1 i_1260 (.A(n_503), .B(n_480), .ZN(n_1368));
   XNOR2_X1 i_1261 (.A(n_1368), .B(n_457), .ZN(n_1369));
   INV_X1 i_1262 (.A(n_1369), .ZN(n_1370));
   OR3_X1 i_1263 (.A1(n_1372), .A2(n_1373), .A3(n_1374), .ZN(n_1371));
   NOR2_X1 i_1264 (.A1(n_480), .A2(n_503), .ZN(n_1372));
   NOR2_X1 i_1265 (.A1(n_457), .A2(n_503), .ZN(n_1373));
   NOR2_X1 i_1266 (.A1(n_457), .A2(n_480), .ZN(n_1374));
   XNOR2_X1 i_1267 (.A(n_434), .B(n_411), .ZN(n_1375));
   XNOR2_X1 i_1268 (.A(n_1375), .B(n_388), .ZN(n_1376));
   INV_X1 i_1269 (.A(n_1376), .ZN(n_1377));
   OR3_X1 i_1270 (.A1(n_1379), .A2(n_1380), .A3(n_1381), .ZN(n_1378));
   NOR2_X1 i_1271 (.A1(n_411), .A2(n_434), .ZN(n_1379));
   NOR2_X1 i_1272 (.A1(n_388), .A2(n_434), .ZN(n_1380));
   NOR2_X1 i_1273 (.A1(n_388), .A2(n_411), .ZN(n_1381));
   XNOR2_X1 i_1274 (.A(n_365), .B(n_342), .ZN(n_1382));
   XNOR2_X1 i_1275 (.A(n_1382), .B(n_319), .ZN(n_1383));
   INV_X1 i_1276 (.A(n_1383), .ZN(n_1384));
   OR3_X1 i_1277 (.A1(n_1386), .A2(n_1387), .A3(n_1388), .ZN(n_1385));
   NOR2_X1 i_1278 (.A1(n_342), .A2(n_365), .ZN(n_1386));
   NOR2_X1 i_1279 (.A1(n_319), .A2(n_365), .ZN(n_1387));
   NOR2_X1 i_1280 (.A1(n_319), .A2(n_342), .ZN(n_1388));
   XNOR2_X1 i_1281 (.A(n_296), .B(n_273), .ZN(n_1389));
   XNOR2_X1 i_1282 (.A(n_1389), .B(n_250), .ZN(n_1390));
   INV_X1 i_1283 (.A(n_1390), .ZN(n_1391));
   OR3_X1 i_1284 (.A1(n_1393), .A2(n_1394), .A3(n_1395), .ZN(n_1392));
   NOR2_X1 i_1285 (.A1(n_273), .A2(n_296), .ZN(n_1393));
   NOR2_X1 i_1286 (.A1(n_250), .A2(n_296), .ZN(n_1394));
   NOR2_X1 i_1287 (.A1(n_250), .A2(n_273), .ZN(n_1395));
   XNOR2_X1 i_1288 (.A(n_227), .B(n_204), .ZN(n_1396));
   XNOR2_X1 i_1289 (.A(n_1396), .B(n_181), .ZN(n_1397));
   INV_X1 i_1290 (.A(n_1397), .ZN(n_1398));
   OR3_X1 i_1291 (.A1(n_1400), .A2(n_1401), .A3(n_1402), .ZN(n_1399));
   NOR2_X1 i_1292 (.A1(n_204), .A2(n_227), .ZN(n_1400));
   NOR2_X1 i_1293 (.A1(n_181), .A2(n_227), .ZN(n_1401));
   NOR2_X1 i_1294 (.A1(n_181), .A2(n_204), .ZN(n_1402));
   XNOR2_X1 i_1295 (.A(n_158), .B(n_135), .ZN(n_1403));
   XNOR2_X1 i_1296 (.A(n_1403), .B(n_112), .ZN(n_1404));
   INV_X1 i_1297 (.A(n_1404), .ZN(n_1405));
   OR3_X1 i_1298 (.A1(n_1407), .A2(n_1408), .A3(n_1409), .ZN(n_1406));
   NOR2_X1 i_1299 (.A1(n_135), .A2(n_158), .ZN(n_1407));
   NOR2_X1 i_1300 (.A1(n_112), .A2(n_158), .ZN(n_1408));
   NOR2_X1 i_1301 (.A1(n_112), .A2(n_135), .ZN(n_1409));
   XNOR2_X1 i_1302 (.A(n_89), .B(n_66), .ZN(n_1410));
   XNOR2_X1 i_1303 (.A(n_1410), .B(n_43), .ZN(n_1411));
   INV_X1 i_1304 (.A(n_1411), .ZN(n_1412));
   OR3_X1 i_1305 (.A1(n_1414), .A2(n_1415), .A3(n_1416), .ZN(n_1413));
   NOR2_X1 i_1306 (.A1(n_66), .A2(n_89), .ZN(n_1414));
   NOR2_X1 i_1307 (.A1(n_43), .A2(n_89), .ZN(n_1415));
   NOR2_X1 i_1308 (.A1(n_43), .A2(n_66), .ZN(n_1416));
   XNOR2_X1 i_1309 (.A(n_20), .B(n_1340), .ZN(n_1417));
   XNOR2_X1 i_1310 (.A(n_1417), .B(n_1333), .ZN(n_1418));
   INV_X1 i_1311 (.A(n_1418), .ZN(n_1419));
   NAND3_X1 i_1312 (.A1(n_1421), .A2(n_1423), .A3(n_1424), .ZN(n_1420));
   NAND2_X1 i_1313 (.A1(n_1340), .A2(n_1422), .ZN(n_1421));
   INV_X1 i_1314 (.A(n_20), .ZN(n_1422));
   NAND2_X1 i_1315 (.A1(n_1333), .A2(n_1422), .ZN(n_1423));
   NAND2_X1 i_1316 (.A1(n_1333), .A2(n_1340), .ZN(n_1424));
   FA_X1 i_1317 (.A(n_1326), .B(n_1319), .CI(n_1312), .CO(n_1426), .S(n_1425));
   FA_X1 i_1318 (.A(n_1305), .B(n_1298), .CI(n_1347), .CO(n_1428), .S(n_1427));
   FA_X1 i_1319 (.A(n_1345), .B(n_1412), .CI(n_1405), .CO(n_1430), .S(n_1429));
   FA_X1 i_1320 (.A(n_1398), .B(n_1391), .CI(n_1384), .CO(n_1432), .S(n_1431));
   FA_X1 i_1321 (.A(n_1377), .B(n_1370), .CI(n_1427), .CO(n_1434), .S(n_1433));
   FA_X1 i_1322 (.A(n_1425), .B(n_1419), .CI(n_1353), .CO(n_1436), .S(n_1435));
   FA_X1 i_1323 (.A(n_1351), .B(n_1349), .CI(n_1355), .CO(n_1438), .S(n_1437));
   FA_X1 i_1324 (.A(n_1433), .B(n_1431), .CI(n_1429), .CO(n_1440), .S(n_1439));
   FA_X1 i_1325 (.A(n_1357), .B(n_1437), .CI(n_1435), .CO(n_1442), .S(n_1441));
   FA_X1 i_1326 (.A(n_1359), .B(n_1361), .CI(n_1439), .CO(n_1444), .S(n_1443));
   FA_X1 i_1327 (.A(n_1363), .B(n_1441), .CI(n_1443), .CO(n_1446), .S(n_1445));
   HA_X1 i_1328 (.A(n_1365), .B(n_1445), .CO(n_1448), .S(n_1447));
   XNOR2_X1 i_1329 (.A(n_527), .B(n_504), .ZN(n_1449));
   XNOR2_X1 i_1330 (.A(n_1449), .B(n_481), .ZN(n_1450));
   INV_X1 i_1331 (.A(n_1450), .ZN(n_1451));
   OR3_X1 i_1332 (.A1(n_1453), .A2(n_1454), .A3(n_1455), .ZN(n_1452));
   NOR2_X1 i_1333 (.A1(n_504), .A2(n_527), .ZN(n_1453));
   NOR2_X1 i_1334 (.A1(n_481), .A2(n_527), .ZN(n_1454));
   NOR2_X1 i_1335 (.A1(n_481), .A2(n_504), .ZN(n_1455));
   XNOR2_X1 i_1336 (.A(n_458), .B(n_435), .ZN(n_1456));
   XNOR2_X1 i_1337 (.A(n_1456), .B(n_412), .ZN(n_1457));
   INV_X1 i_1338 (.A(n_1457), .ZN(n_1458));
   OR3_X1 i_1339 (.A1(n_1460), .A2(n_1461), .A3(n_1462), .ZN(n_1459));
   NOR2_X1 i_1340 (.A1(n_435), .A2(n_458), .ZN(n_1460));
   NOR2_X1 i_1341 (.A1(n_412), .A2(n_458), .ZN(n_1461));
   NOR2_X1 i_1342 (.A1(n_412), .A2(n_435), .ZN(n_1462));
   XNOR2_X1 i_1343 (.A(n_389), .B(n_366), .ZN(n_1463));
   XNOR2_X1 i_1344 (.A(n_1463), .B(n_343), .ZN(n_1464));
   INV_X1 i_1345 (.A(n_1464), .ZN(n_1465));
   OR3_X1 i_1346 (.A1(n_1467), .A2(n_1468), .A3(n_1469), .ZN(n_1466));
   NOR2_X1 i_1347 (.A1(n_366), .A2(n_389), .ZN(n_1467));
   NOR2_X1 i_1348 (.A1(n_343), .A2(n_389), .ZN(n_1468));
   NOR2_X1 i_1349 (.A1(n_343), .A2(n_366), .ZN(n_1469));
   XNOR2_X1 i_1350 (.A(n_320), .B(n_297), .ZN(n_1470));
   XNOR2_X1 i_1351 (.A(n_1470), .B(n_274), .ZN(n_1471));
   INV_X1 i_1352 (.A(n_1471), .ZN(n_1472));
   OR3_X1 i_1353 (.A1(n_1474), .A2(n_1475), .A3(n_1476), .ZN(n_1473));
   NOR2_X1 i_1354 (.A1(n_297), .A2(n_320), .ZN(n_1474));
   NOR2_X1 i_1355 (.A1(n_274), .A2(n_320), .ZN(n_1475));
   NOR2_X1 i_1356 (.A1(n_274), .A2(n_297), .ZN(n_1476));
   XNOR2_X1 i_1357 (.A(n_251), .B(n_228), .ZN(n_1477));
   XNOR2_X1 i_1358 (.A(n_1477), .B(n_205), .ZN(n_1478));
   INV_X1 i_1359 (.A(n_1478), .ZN(n_1479));
   OR3_X1 i_1360 (.A1(n_1481), .A2(n_1482), .A3(n_1483), .ZN(n_1480));
   NOR2_X1 i_1361 (.A1(n_228), .A2(n_251), .ZN(n_1481));
   NOR2_X1 i_1362 (.A1(n_205), .A2(n_251), .ZN(n_1482));
   NOR2_X1 i_1363 (.A1(n_205), .A2(n_228), .ZN(n_1483));
   XNOR2_X1 i_1364 (.A(n_182), .B(n_159), .ZN(n_1484));
   XNOR2_X1 i_1365 (.A(n_1484), .B(n_136), .ZN(n_1485));
   INV_X1 i_1366 (.A(n_1485), .ZN(n_1486));
   OR3_X1 i_1367 (.A1(n_1488), .A2(n_1489), .A3(n_1490), .ZN(n_1487));
   NOR2_X1 i_1368 (.A1(n_159), .A2(n_182), .ZN(n_1488));
   NOR2_X1 i_1369 (.A1(n_136), .A2(n_182), .ZN(n_1489));
   NOR2_X1 i_1370 (.A1(n_136), .A2(n_159), .ZN(n_1490));
   XNOR2_X1 i_1371 (.A(n_113), .B(n_90), .ZN(n_1491));
   XNOR2_X1 i_1372 (.A(n_1491), .B(n_67), .ZN(n_1492));
   INV_X1 i_1373 (.A(n_1492), .ZN(n_1493));
   OR3_X1 i_1374 (.A1(n_1495), .A2(n_1496), .A3(n_1497), .ZN(n_1494));
   NOR2_X1 i_1375 (.A1(n_90), .A2(n_113), .ZN(n_1495));
   NOR2_X1 i_1376 (.A1(n_67), .A2(n_113), .ZN(n_1496));
   NOR2_X1 i_1377 (.A1(n_67), .A2(n_90), .ZN(n_1497));
   XNOR2_X1 i_1378 (.A(n_44), .B(n_21), .ZN(n_1498));
   XNOR2_X1 i_1379 (.A(n_1498), .B(n_1413), .ZN(n_1499));
   NAND3_X1 i_1380 (.A1(n_1501), .A2(n_1502), .A3(n_1504), .ZN(n_1500));
   OR2_X1 i_1381 (.A1(n_21), .A2(n_44), .ZN(n_1501));
   NAND2_X1 i_1382 (.A1(n_1413), .A2(n_1503), .ZN(n_1502));
   INV_X1 i_1383 (.A(n_44), .ZN(n_1503));
   NAND2_X1 i_1384 (.A1(n_1413), .A2(n_1505), .ZN(n_1504));
   INV_X1 i_1385 (.A(n_21), .ZN(n_1505));
   FA_X1 i_1386 (.A(n_1406), .B(n_1399), .CI(n_1392), .CO(n_1507), .S(n_1506));
   FA_X1 i_1387 (.A(n_1385), .B(n_1378), .CI(n_1371), .CO(n_1509), .S(n_1508));
   FA_X1 i_1388 (.A(n_1426), .B(n_1420), .CI(n_1499), .CO(n_1511), .S(n_1510));
   FA_X1 i_1389 (.A(n_1493), .B(n_1486), .CI(n_1479), .CO(n_1513), .S(n_1512));
   FA_X1 i_1390 (.A(n_1472), .B(n_1465), .CI(n_1458), .CO(n_1515), .S(n_1514));
   FA_X1 i_1391 (.A(n_1451), .B(n_1428), .CI(n_1508), .CO(n_1517), .S(n_1516));
   FA_X1 i_1392 (.A(n_1506), .B(n_1432), .CI(n_1430), .CO(n_1519), .S(n_1518));
   FA_X1 i_1393 (.A(n_1510), .B(n_1436), .CI(n_1434), .CO(n_1521), .S(n_1520));
   FA_X1 i_1394 (.A(n_1514), .B(n_1512), .CI(n_1516), .CO(n_1523), .S(n_1522));
   FA_X1 i_1395 (.A(n_1438), .B(n_1518), .CI(n_1440), .CO(n_1525), .S(n_1524));
   FA_X1 i_1396 (.A(n_1520), .B(n_1442), .CI(n_1522), .CO(n_1527), .S(n_1526));
   FA_X1 i_1397 (.A(n_1524), .B(n_1444), .CI(n_1526), .CO(n_1529), .S(n_1528));
   HA_X1 i_1398 (.A(n_1446), .B(n_1528), .CO(n_1531), .S(n_1530));
   XNOR2_X1 i_1399 (.A(n_551), .B(n_528), .ZN(n_1532));
   XNOR2_X1 i_1400 (.A(n_1532), .B(n_505), .ZN(n_1533));
   INV_X1 i_1401 (.A(n_1533), .ZN(n_1534));
   OR3_X1 i_1402 (.A1(n_1536), .A2(n_1537), .A3(n_1538), .ZN(n_1535));
   NOR2_X1 i_1403 (.A1(n_528), .A2(n_551), .ZN(n_1536));
   NOR2_X1 i_1404 (.A1(n_505), .A2(n_551), .ZN(n_1537));
   NOR2_X1 i_1405 (.A1(n_505), .A2(n_528), .ZN(n_1538));
   XNOR2_X1 i_1406 (.A(n_482), .B(n_459), .ZN(n_1539));
   XNOR2_X1 i_1407 (.A(n_1539), .B(n_436), .ZN(n_1540));
   INV_X1 i_1408 (.A(n_1540), .ZN(n_1541));
   OR3_X1 i_1409 (.A1(n_1543), .A2(n_1544), .A3(n_1545), .ZN(n_1542));
   NOR2_X1 i_1410 (.A1(n_459), .A2(n_482), .ZN(n_1543));
   NOR2_X1 i_1411 (.A1(n_436), .A2(n_482), .ZN(n_1544));
   NOR2_X1 i_1412 (.A1(n_436), .A2(n_459), .ZN(n_1545));
   XNOR2_X1 i_1413 (.A(n_413), .B(n_390), .ZN(n_1546));
   XNOR2_X1 i_1414 (.A(n_1546), .B(n_367), .ZN(n_1547));
   INV_X1 i_1415 (.A(n_1547), .ZN(n_1548));
   OR3_X1 i_1416 (.A1(n_1550), .A2(n_1551), .A3(n_1552), .ZN(n_1549));
   NOR2_X1 i_1417 (.A1(n_390), .A2(n_413), .ZN(n_1550));
   NOR2_X1 i_1418 (.A1(n_367), .A2(n_413), .ZN(n_1551));
   NOR2_X1 i_1419 (.A1(n_367), .A2(n_390), .ZN(n_1552));
   XNOR2_X1 i_1420 (.A(n_344), .B(n_321), .ZN(n_1553));
   XNOR2_X1 i_1421 (.A(n_1553), .B(n_298), .ZN(n_1554));
   INV_X1 i_1422 (.A(n_1554), .ZN(n_1555));
   OR3_X1 i_1423 (.A1(n_1557), .A2(n_1558), .A3(n_1559), .ZN(n_1556));
   NOR2_X1 i_1424 (.A1(n_321), .A2(n_344), .ZN(n_1557));
   NOR2_X1 i_1425 (.A1(n_298), .A2(n_344), .ZN(n_1558));
   NOR2_X1 i_1426 (.A1(n_298), .A2(n_321), .ZN(n_1559));
   XNOR2_X1 i_1427 (.A(n_275), .B(n_252), .ZN(n_1560));
   XNOR2_X1 i_1428 (.A(n_1560), .B(n_229), .ZN(n_1561));
   INV_X1 i_1429 (.A(n_1561), .ZN(n_1562));
   OR3_X1 i_1430 (.A1(n_1564), .A2(n_1565), .A3(n_1566), .ZN(n_1563));
   NOR2_X1 i_1431 (.A1(n_252), .A2(n_275), .ZN(n_1564));
   NOR2_X1 i_1432 (.A1(n_229), .A2(n_275), .ZN(n_1565));
   NOR2_X1 i_1433 (.A1(n_229), .A2(n_252), .ZN(n_1566));
   XNOR2_X1 i_1434 (.A(n_206), .B(n_183), .ZN(n_1567));
   XNOR2_X1 i_1435 (.A(n_1567), .B(n_160), .ZN(n_1568));
   INV_X1 i_1436 (.A(n_1568), .ZN(n_1569));
   OR3_X1 i_1437 (.A1(n_1571), .A2(n_1572), .A3(n_1573), .ZN(n_1570));
   NOR2_X1 i_1438 (.A1(n_183), .A2(n_206), .ZN(n_1571));
   NOR2_X1 i_1439 (.A1(n_160), .A2(n_206), .ZN(n_1572));
   NOR2_X1 i_1440 (.A1(n_160), .A2(n_183), .ZN(n_1573));
   XNOR2_X1 i_1441 (.A(n_137), .B(n_114), .ZN(n_1574));
   XNOR2_X1 i_1442 (.A(n_1574), .B(n_91), .ZN(n_1575));
   INV_X1 i_1443 (.A(n_1575), .ZN(n_1576));
   OR3_X1 i_1444 (.A1(n_1578), .A2(n_1579), .A3(n_1580), .ZN(n_1577));
   NOR2_X1 i_1445 (.A1(n_114), .A2(n_137), .ZN(n_1578));
   NOR2_X1 i_1446 (.A1(n_91), .A2(n_137), .ZN(n_1579));
   NOR2_X1 i_1447 (.A1(n_91), .A2(n_114), .ZN(n_1580));
   XNOR2_X1 i_1448 (.A(n_68), .B(n_45), .ZN(n_1581));
   XNOR2_X1 i_1449 (.A(n_1581), .B(n_22), .ZN(n_1582));
   INV_X1 i_1450 (.A(n_1582), .ZN(n_1583));
   OR3_X1 i_1451 (.A1(n_1585), .A2(n_1586), .A3(n_1587), .ZN(n_1584));
   NOR2_X1 i_1452 (.A1(n_45), .A2(n_68), .ZN(n_1585));
   NOR2_X1 i_1453 (.A1(n_22), .A2(n_68), .ZN(n_1586));
   NOR2_X1 i_1454 (.A1(n_22), .A2(n_45), .ZN(n_1587));
   FA_X1 i_1455 (.A(n_1494), .B(n_1487), .CI(n_1480), .CO(n_1589), .S(n_1588));
   FA_X1 i_1456 (.A(n_1473), .B(n_1466), .CI(n_1459), .CO(n_1591), .S(n_1590));
   FA_X1 i_1457 (.A(n_1452), .B(n_1509), .CI(n_1507), .CO(n_1593), .S(n_1592));
   FA_X1 i_1458 (.A(n_1500), .B(n_1583), .CI(n_1576), .CO(n_1595), .S(n_1594));
   FA_X1 i_1459 (.A(n_1569), .B(n_1562), .CI(n_1555), .CO(n_1597), .S(n_1596));
   FA_X1 i_1460 (.A(n_1548), .B(n_1541), .CI(n_1534), .CO(n_1599), .S(n_1598));
   FA_X1 i_1461 (.A(n_1590), .B(n_1588), .CI(n_1515), .CO(n_1601), .S(n_1600));
   FA_X1 i_1462 (.A(n_1513), .B(n_1511), .CI(n_1592), .CO(n_1603), .S(n_1602));
   FA_X1 i_1463 (.A(n_1519), .B(n_1517), .CI(n_1598), .CO(n_1605), .S(n_1604));
   FA_X1 i_1464 (.A(n_1596), .B(n_1594), .CI(n_1521), .CO(n_1607), .S(n_1606));
   FA_X1 i_1465 (.A(n_1602), .B(n_1600), .CI(n_1523), .CO(n_1609), .S(n_1608));
   FA_X1 i_1466 (.A(n_1604), .B(n_1525), .CI(n_1606), .CO(n_1611), .S(n_1610));
   FA_X1 i_1467 (.A(n_1608), .B(n_1527), .CI(n_1610), .CO(n_1613), .S(n_1612));
   HA_X1 i_1468 (.A(n_1529), .B(n_1612), .CO(n_1615), .S(n_1614));
   XNOR2_X1 i_1469 (.A(n_552), .B(n_529), .ZN(n_1616));
   XNOR2_X1 i_1470 (.A(n_1616), .B(n_506), .ZN(n_1617));
   INV_X1 i_1471 (.A(n_1617), .ZN(n_1618));
   OR3_X1 i_1472 (.A1(n_1620), .A2(n_1621), .A3(n_1622), .ZN(n_1619));
   NOR2_X1 i_1473 (.A1(n_529), .A2(n_552), .ZN(n_1620));
   NOR2_X1 i_1474 (.A1(n_506), .A2(n_552), .ZN(n_1621));
   NOR2_X1 i_1475 (.A1(n_506), .A2(n_529), .ZN(n_1622));
   XNOR2_X1 i_1476 (.A(n_483), .B(n_460), .ZN(n_1623));
   XNOR2_X1 i_1477 (.A(n_1623), .B(n_437), .ZN(n_1624));
   INV_X1 i_1478 (.A(n_1624), .ZN(n_1625));
   OR3_X1 i_1479 (.A1(n_1627), .A2(n_1628), .A3(n_1629), .ZN(n_1626));
   NOR2_X1 i_1480 (.A1(n_460), .A2(n_483), .ZN(n_1627));
   NOR2_X1 i_1481 (.A1(n_437), .A2(n_483), .ZN(n_1628));
   NOR2_X1 i_1482 (.A1(n_437), .A2(n_460), .ZN(n_1629));
   XNOR2_X1 i_1483 (.A(n_414), .B(n_391), .ZN(n_1630));
   XNOR2_X1 i_1484 (.A(n_1630), .B(n_368), .ZN(n_1631));
   INV_X1 i_1485 (.A(n_1631), .ZN(n_1632));
   OR3_X1 i_1486 (.A1(n_1634), .A2(n_1635), .A3(n_1636), .ZN(n_1633));
   NOR2_X1 i_1487 (.A1(n_391), .A2(n_414), .ZN(n_1634));
   NOR2_X1 i_1488 (.A1(n_368), .A2(n_414), .ZN(n_1635));
   NOR2_X1 i_1489 (.A1(n_368), .A2(n_391), .ZN(n_1636));
   XNOR2_X1 i_1490 (.A(n_345), .B(n_322), .ZN(n_1637));
   XNOR2_X1 i_1491 (.A(n_1637), .B(n_299), .ZN(n_1638));
   INV_X1 i_1492 (.A(n_1638), .ZN(n_1639));
   OR3_X1 i_1493 (.A1(n_1641), .A2(n_1642), .A3(n_1643), .ZN(n_1640));
   NOR2_X1 i_1494 (.A1(n_322), .A2(n_345), .ZN(n_1641));
   NOR2_X1 i_1495 (.A1(n_299), .A2(n_345), .ZN(n_1642));
   NOR2_X1 i_1496 (.A1(n_299), .A2(n_322), .ZN(n_1643));
   XNOR2_X1 i_1497 (.A(n_276), .B(n_253), .ZN(n_1644));
   XNOR2_X1 i_1498 (.A(n_1644), .B(n_230), .ZN(n_1645));
   INV_X1 i_1499 (.A(n_1645), .ZN(n_1646));
   OR3_X1 i_1500 (.A1(n_1648), .A2(n_1649), .A3(n_1650), .ZN(n_1647));
   NOR2_X1 i_1501 (.A1(n_253), .A2(n_276), .ZN(n_1648));
   NOR2_X1 i_1502 (.A1(n_230), .A2(n_276), .ZN(n_1649));
   NOR2_X1 i_1503 (.A1(n_230), .A2(n_253), .ZN(n_1650));
   XNOR2_X1 i_1504 (.A(n_207), .B(n_184), .ZN(n_1651));
   XNOR2_X1 i_1505 (.A(n_1651), .B(n_161), .ZN(n_1652));
   INV_X1 i_1506 (.A(n_1652), .ZN(n_1653));
   OR3_X1 i_1507 (.A1(n_1655), .A2(n_1656), .A3(n_1657), .ZN(n_1654));
   NOR2_X1 i_1508 (.A1(n_184), .A2(n_207), .ZN(n_1655));
   NOR2_X1 i_1509 (.A1(n_161), .A2(n_207), .ZN(n_1656));
   NOR2_X1 i_1510 (.A1(n_161), .A2(n_184), .ZN(n_1657));
   XNOR2_X1 i_1511 (.A(n_138), .B(n_115), .ZN(n_1658));
   XNOR2_X1 i_1512 (.A(n_1658), .B(n_92), .ZN(n_1659));
   INV_X1 i_1513 (.A(n_1659), .ZN(n_1660));
   OR3_X1 i_1514 (.A1(n_1662), .A2(n_1663), .A3(n_1664), .ZN(n_1661));
   NOR2_X1 i_1515 (.A1(n_115), .A2(n_138), .ZN(n_1662));
   NOR2_X1 i_1516 (.A1(n_92), .A2(n_138), .ZN(n_1663));
   NOR2_X1 i_1517 (.A1(n_92), .A2(n_115), .ZN(n_1664));
   XNOR2_X1 i_1518 (.A(n_69), .B(n_46), .ZN(n_1665));
   XNOR2_X1 i_1519 (.A(n_1665), .B(n_1584), .ZN(n_1666));
   NAND3_X1 i_1520 (.A1(n_1668), .A2(n_1669), .A3(n_1671), .ZN(n_1667));
   OR2_X1 i_1521 (.A1(n_46), .A2(n_69), .ZN(n_1668));
   NAND2_X1 i_1522 (.A1(n_1584), .A2(n_1670), .ZN(n_1669));
   INV_X1 i_1523 (.A(n_69), .ZN(n_1670));
   NAND2_X1 i_1524 (.A1(n_1584), .A2(n_1672), .ZN(n_1671));
   INV_X1 i_1525 (.A(n_46), .ZN(n_1672));
   FA_X1 i_1526 (.A(n_1577), .B(n_1570), .CI(n_1563), .CO(n_1674), .S(n_1673));
   FA_X1 i_1527 (.A(n_1556), .B(n_1549), .CI(n_1542), .CO(n_1676), .S(n_1675));
   FA_X1 i_1528 (.A(n_1535), .B(n_1591), .CI(n_1589), .CO(n_1678), .S(n_1677));
   FA_X1 i_1529 (.A(n_1666), .B(n_1660), .CI(n_1653), .CO(n_1680), .S(n_1679));
   FA_X1 i_1530 (.A(n_1646), .B(n_1639), .CI(n_1632), .CO(n_1682), .S(n_1681));
   FA_X1 i_1531 (.A(n_1625), .B(n_1618), .CI(n_1593), .CO(n_1684), .S(n_1683));
   FA_X1 i_1532 (.A(n_1675), .B(n_1673), .CI(n_1599), .CO(n_1686), .S(n_1685));
   FA_X1 i_1533 (.A(n_1597), .B(n_1595), .CI(n_1677), .CO(n_1688), .S(n_1687));
   FA_X1 i_1534 (.A(n_1601), .B(n_1683), .CI(n_1681), .CO(n_1690), .S(n_1689));
   FA_X1 i_1535 (.A(n_1679), .B(n_1603), .CI(n_1687), .CO(n_1692), .S(n_1691));
   FA_X1 i_1536 (.A(n_1685), .B(n_1605), .CI(n_1607), .CO(n_1694), .S(n_1693));
   FA_X1 i_1537 (.A(n_1609), .B(n_1689), .CI(n_1691), .CO(n_1696), .S(n_1695));
   FA_X1 i_1538 (.A(n_1693), .B(n_1611), .CI(n_1695), .CO(n_1698), .S(n_1697));
   HA_X1 i_1539 (.A(n_1613), .B(n_1697), .CO(n_1700), .S(n_1699));
   XNOR2_X1 i_1540 (.A(n_553), .B(n_530), .ZN(n_1701));
   XNOR2_X1 i_1541 (.A(n_1701), .B(n_507), .ZN(n_1702));
   INV_X1 i_1542 (.A(n_1702), .ZN(n_1703));
   OR3_X1 i_1543 (.A1(n_1705), .A2(n_1706), .A3(n_1707), .ZN(n_1704));
   NOR2_X1 i_1544 (.A1(n_530), .A2(n_553), .ZN(n_1705));
   NOR2_X1 i_1545 (.A1(n_507), .A2(n_553), .ZN(n_1706));
   NOR2_X1 i_1546 (.A1(n_507), .A2(n_530), .ZN(n_1707));
   XNOR2_X1 i_1547 (.A(n_484), .B(n_461), .ZN(n_1708));
   XNOR2_X1 i_1548 (.A(n_1708), .B(n_438), .ZN(n_1709));
   INV_X1 i_1549 (.A(n_1709), .ZN(n_1710));
   OR3_X1 i_1550 (.A1(n_1712), .A2(n_1713), .A3(n_1714), .ZN(n_1711));
   NOR2_X1 i_1551 (.A1(n_461), .A2(n_484), .ZN(n_1712));
   NOR2_X1 i_1552 (.A1(n_438), .A2(n_484), .ZN(n_1713));
   NOR2_X1 i_1553 (.A1(n_438), .A2(n_461), .ZN(n_1714));
   XNOR2_X1 i_1554 (.A(n_415), .B(n_392), .ZN(n_1715));
   XNOR2_X1 i_1555 (.A(n_1715), .B(n_369), .ZN(n_1716));
   INV_X1 i_1556 (.A(n_1716), .ZN(n_1717));
   OR3_X1 i_1557 (.A1(n_1719), .A2(n_1720), .A3(n_1721), .ZN(n_1718));
   NOR2_X1 i_1558 (.A1(n_392), .A2(n_415), .ZN(n_1719));
   NOR2_X1 i_1559 (.A1(n_369), .A2(n_415), .ZN(n_1720));
   NOR2_X1 i_1560 (.A1(n_369), .A2(n_392), .ZN(n_1721));
   XNOR2_X1 i_1561 (.A(n_346), .B(n_323), .ZN(n_1722));
   XNOR2_X1 i_1562 (.A(n_1722), .B(n_300), .ZN(n_1723));
   INV_X1 i_1563 (.A(n_1723), .ZN(n_1724));
   OR3_X1 i_1564 (.A1(n_1726), .A2(n_1727), .A3(n_1728), .ZN(n_1725));
   NOR2_X1 i_1565 (.A1(n_323), .A2(n_346), .ZN(n_1726));
   NOR2_X1 i_1566 (.A1(n_300), .A2(n_346), .ZN(n_1727));
   NOR2_X1 i_1567 (.A1(n_300), .A2(n_323), .ZN(n_1728));
   XNOR2_X1 i_1568 (.A(n_277), .B(n_254), .ZN(n_1729));
   XNOR2_X1 i_1569 (.A(n_1729), .B(n_231), .ZN(n_1730));
   INV_X1 i_1570 (.A(n_1730), .ZN(n_1731));
   OR3_X1 i_1571 (.A1(n_1733), .A2(n_1734), .A3(n_1735), .ZN(n_1732));
   NOR2_X1 i_1572 (.A1(n_254), .A2(n_277), .ZN(n_1733));
   NOR2_X1 i_1573 (.A1(n_231), .A2(n_277), .ZN(n_1734));
   NOR2_X1 i_1574 (.A1(n_231), .A2(n_254), .ZN(n_1735));
   XNOR2_X1 i_1575 (.A(n_208), .B(n_185), .ZN(n_1736));
   XNOR2_X1 i_1576 (.A(n_1736), .B(n_162), .ZN(n_1737));
   INV_X1 i_1577 (.A(n_1737), .ZN(n_1738));
   OR3_X1 i_1578 (.A1(n_1740), .A2(n_1741), .A3(n_1742), .ZN(n_1739));
   NOR2_X1 i_1579 (.A1(n_185), .A2(n_208), .ZN(n_1740));
   NOR2_X1 i_1580 (.A1(n_162), .A2(n_208), .ZN(n_1741));
   NOR2_X1 i_1581 (.A1(n_162), .A2(n_185), .ZN(n_1742));
   XNOR2_X1 i_1582 (.A(n_139), .B(n_116), .ZN(n_1743));
   XNOR2_X1 i_1583 (.A(n_1743), .B(n_93), .ZN(n_1744));
   INV_X1 i_1584 (.A(n_1744), .ZN(n_1745));
   OR3_X1 i_1585 (.A1(n_1747), .A2(n_1748), .A3(n_1749), .ZN(n_1746));
   NOR2_X1 i_1586 (.A1(n_116), .A2(n_139), .ZN(n_1747));
   NOR2_X1 i_1587 (.A1(n_93), .A2(n_139), .ZN(n_1748));
   NOR2_X1 i_1588 (.A1(n_93), .A2(n_116), .ZN(n_1749));
   XNOR2_X1 i_1589 (.A(n_70), .B(n_1661), .ZN(n_1750));
   XNOR2_X1 i_1590 (.A(n_1750), .B(n_1654), .ZN(n_1751));
   INV_X1 i_1591 (.A(n_1751), .ZN(n_1752));
   NAND3_X1 i_1592 (.A1(n_1754), .A2(n_1756), .A3(n_1757), .ZN(n_1753));
   NAND2_X1 i_1593 (.A1(n_1661), .A2(n_1755), .ZN(n_1754));
   INV_X1 i_1594 (.A(n_70), .ZN(n_1755));
   NAND2_X1 i_1595 (.A1(n_1654), .A2(n_1755), .ZN(n_1756));
   NAND2_X1 i_1596 (.A1(n_1654), .A2(n_1661), .ZN(n_1757));
   FA_X1 i_1597 (.A(n_1647), .B(n_1640), .CI(n_1633), .CO(n_1759), .S(n_1758));
   FA_X1 i_1598 (.A(n_1626), .B(n_1619), .CI(n_1676), .CO(n_1761), .S(n_1760));
   FA_X1 i_1599 (.A(n_1674), .B(n_1667), .CI(n_1745), .CO(n_1763), .S(n_1762));
   FA_X1 i_1600 (.A(n_1738), .B(n_1731), .CI(n_1724), .CO(n_1765), .S(n_1764));
   FA_X1 i_1601 (.A(n_1717), .B(n_1710), .CI(n_1703), .CO(n_1767), .S(n_1766));
   FA_X1 i_1602 (.A(n_1678), .B(n_1760), .CI(n_1758), .CO(n_1769), .S(n_1768));
   FA_X1 i_1603 (.A(n_1752), .B(n_1682), .CI(n_1680), .CO(n_1771), .S(n_1770));
   FA_X1 i_1604 (.A(n_1684), .B(n_1762), .CI(n_1686), .CO(n_1773), .S(n_1772));
   FA_X1 i_1605 (.A(n_1766), .B(n_1764), .CI(n_1688), .CO(n_1775), .S(n_1774));
   FA_X1 i_1606 (.A(n_1770), .B(n_1768), .CI(n_1690), .CO(n_1777), .S(n_1776));
   FA_X1 i_1607 (.A(n_1772), .B(n_1692), .CI(n_1694), .CO(n_1779), .S(n_1778));
   FA_X1 i_1608 (.A(n_1774), .B(n_1776), .CI(n_1696), .CO(n_1781), .S(n_1780));
   FA_X1 i_1609 (.A(n_1778), .B(n_1780), .CI(n_1698), .CO(n_1783), .S(n_1782));
   XNOR2_X1 i_1610 (.A(n_554), .B(n_531), .ZN(n_1784));
   XNOR2_X1 i_1611 (.A(n_1784), .B(n_508), .ZN(n_1785));
   INV_X1 i_1612 (.A(n_1785), .ZN(n_1786));
   OR3_X1 i_1613 (.A1(n_1788), .A2(n_1789), .A3(n_1790), .ZN(n_1787));
   NOR2_X1 i_1614 (.A1(n_531), .A2(n_554), .ZN(n_1788));
   NOR2_X1 i_1615 (.A1(n_508), .A2(n_554), .ZN(n_1789));
   NOR2_X1 i_1616 (.A1(n_508), .A2(n_531), .ZN(n_1790));
   XNOR2_X1 i_1617 (.A(n_485), .B(n_462), .ZN(n_1791));
   XNOR2_X1 i_1618 (.A(n_1791), .B(n_439), .ZN(n_1792));
   INV_X1 i_1619 (.A(n_1792), .ZN(n_1793));
   OR3_X1 i_1620 (.A1(n_1795), .A2(n_1796), .A3(n_1797), .ZN(n_1794));
   NOR2_X1 i_1621 (.A1(n_462), .A2(n_485), .ZN(n_1795));
   NOR2_X1 i_1622 (.A1(n_439), .A2(n_485), .ZN(n_1796));
   NOR2_X1 i_1623 (.A1(n_439), .A2(n_462), .ZN(n_1797));
   XNOR2_X1 i_1624 (.A(n_416), .B(n_393), .ZN(n_1798));
   XNOR2_X1 i_1625 (.A(n_1798), .B(n_370), .ZN(n_1799));
   INV_X1 i_1626 (.A(n_1799), .ZN(n_1800));
   OR3_X1 i_1627 (.A1(n_1802), .A2(n_1803), .A3(n_1804), .ZN(n_1801));
   NOR2_X1 i_1628 (.A1(n_393), .A2(n_416), .ZN(n_1802));
   NOR2_X1 i_1629 (.A1(n_370), .A2(n_416), .ZN(n_1803));
   NOR2_X1 i_1630 (.A1(n_370), .A2(n_393), .ZN(n_1804));
   XNOR2_X1 i_1631 (.A(n_347), .B(n_324), .ZN(n_1805));
   XNOR2_X1 i_1632 (.A(n_1805), .B(n_301), .ZN(n_1806));
   INV_X1 i_1633 (.A(n_1806), .ZN(n_1807));
   OR3_X1 i_1634 (.A1(n_1809), .A2(n_1810), .A3(n_1811), .ZN(n_1808));
   NOR2_X1 i_1635 (.A1(n_324), .A2(n_347), .ZN(n_1809));
   NOR2_X1 i_1636 (.A1(n_301), .A2(n_347), .ZN(n_1810));
   NOR2_X1 i_1637 (.A1(n_301), .A2(n_324), .ZN(n_1811));
   XNOR2_X1 i_1638 (.A(n_278), .B(n_255), .ZN(n_1812));
   XNOR2_X1 i_1639 (.A(n_1812), .B(n_232), .ZN(n_1813));
   INV_X1 i_1640 (.A(n_1813), .ZN(n_1814));
   OR3_X1 i_1641 (.A1(n_1816), .A2(n_1817), .A3(n_1818), .ZN(n_1815));
   NOR2_X1 i_1642 (.A1(n_255), .A2(n_278), .ZN(n_1816));
   NOR2_X1 i_1643 (.A1(n_232), .A2(n_278), .ZN(n_1817));
   NOR2_X1 i_1644 (.A1(n_232), .A2(n_255), .ZN(n_1818));
   XNOR2_X1 i_1645 (.A(n_209), .B(n_186), .ZN(n_1819));
   XNOR2_X1 i_1646 (.A(n_1819), .B(n_163), .ZN(n_1820));
   INV_X1 i_1647 (.A(n_1820), .ZN(n_1821));
   OR3_X1 i_1648 (.A1(n_1823), .A2(n_1824), .A3(n_1825), .ZN(n_1822));
   NOR2_X1 i_1649 (.A1(n_186), .A2(n_209), .ZN(n_1823));
   NOR2_X1 i_1650 (.A1(n_163), .A2(n_209), .ZN(n_1824));
   NOR2_X1 i_1651 (.A1(n_163), .A2(n_186), .ZN(n_1825));
   XNOR2_X1 i_1652 (.A(n_140), .B(n_117), .ZN(n_1826));
   XNOR2_X1 i_1653 (.A(n_1826), .B(n_94), .ZN(n_1827));
   INV_X1 i_1654 (.A(n_1827), .ZN(n_1828));
   OR3_X1 i_1655 (.A1(n_1830), .A2(n_1831), .A3(n_1832), .ZN(n_1829));
   NOR2_X1 i_1656 (.A1(n_117), .A2(n_140), .ZN(n_1830));
   NOR2_X1 i_1657 (.A1(n_94), .A2(n_140), .ZN(n_1831));
   NOR2_X1 i_1658 (.A1(n_94), .A2(n_117), .ZN(n_1832));
   FA_X1 i_1659 (.A(n_1746), .B(n_1739), .CI(n_1732), .CO(n_1834), .S(n_1833));
   FA_X1 i_1660 (.A(n_1725), .B(n_1718), .CI(n_1711), .CO(n_1836), .S(n_1835));
   FA_X1 i_1661 (.A(n_1704), .B(n_1759), .CI(n_1753), .CO(n_1838), .S(n_1837));
   FA_X1 i_1662 (.A(n_1828), .B(n_1821), .CI(n_1814), .CO(n_1840), .S(n_1839));
   FA_X1 i_1663 (.A(n_1807), .B(n_1800), .CI(n_1793), .CO(n_1842), .S(n_1841));
   FA_X1 i_1664 (.A(n_1786), .B(n_1761), .CI(n_1835), .CO(n_1844), .S(n_1843));
   FA_X1 i_1665 (.A(n_1833), .B(n_1767), .CI(n_1765), .CO(n_1846), .S(n_1845));
   FA_X1 i_1666 (.A(n_1763), .B(n_1837), .CI(n_1771), .CO(n_1848), .S(n_1847));
   FA_X1 i_1667 (.A(n_1769), .B(n_1841), .CI(n_1839), .CO(n_1850), .S(n_1849));
   FA_X1 i_1668 (.A(n_1843), .B(n_1773), .CI(n_1845), .CO(n_1852), .S(n_1851));
   FA_X1 i_1669 (.A(n_1775), .B(n_1847), .CI(n_1777), .CO(n_1854), .S(n_1853));
   FA_X1 i_1670 (.A(n_1849), .B(n_1851), .CI(n_1779), .CO(n_1856), .S(n_1855));
   FA_X1 i_1671 (.A(n_1853), .B(n_1781), .CI(n_1855), .CO(n_1858), .S(n_1857));
   XNOR2_X1 i_1672 (.A(n_555), .B(n_532), .ZN(n_1859));
   XNOR2_X1 i_1673 (.A(n_1859), .B(n_509), .ZN(n_1860));
   INV_X1 i_1674 (.A(n_1860), .ZN(n_1861));
   OR3_X1 i_1675 (.A1(n_1863), .A2(n_1864), .A3(n_1865), .ZN(n_1862));
   NOR2_X1 i_1676 (.A1(n_532), .A2(n_555), .ZN(n_1863));
   NOR2_X1 i_1677 (.A1(n_509), .A2(n_555), .ZN(n_1864));
   NOR2_X1 i_1678 (.A1(n_509), .A2(n_532), .ZN(n_1865));
   XNOR2_X1 i_1679 (.A(n_486), .B(n_463), .ZN(n_1866));
   XNOR2_X1 i_1680 (.A(n_1866), .B(n_440), .ZN(n_1867));
   INV_X1 i_1681 (.A(n_1867), .ZN(n_1868));
   OR3_X1 i_1682 (.A1(n_1870), .A2(n_1871), .A3(n_1872), .ZN(n_1869));
   NOR2_X1 i_1683 (.A1(n_463), .A2(n_486), .ZN(n_1870));
   NOR2_X1 i_1684 (.A1(n_440), .A2(n_486), .ZN(n_1871));
   NOR2_X1 i_1685 (.A1(n_440), .A2(n_463), .ZN(n_1872));
   XNOR2_X1 i_1686 (.A(n_417), .B(n_394), .ZN(n_1873));
   XNOR2_X1 i_1687 (.A(n_1873), .B(n_371), .ZN(n_1874));
   INV_X1 i_1688 (.A(n_1874), .ZN(n_1875));
   OR3_X1 i_1689 (.A1(n_1877), .A2(n_1878), .A3(n_1879), .ZN(n_1876));
   NOR2_X1 i_1690 (.A1(n_394), .A2(n_417), .ZN(n_1877));
   NOR2_X1 i_1691 (.A1(n_371), .A2(n_417), .ZN(n_1878));
   NOR2_X1 i_1692 (.A1(n_371), .A2(n_394), .ZN(n_1879));
   XNOR2_X1 i_1693 (.A(n_348), .B(n_325), .ZN(n_1880));
   XNOR2_X1 i_1694 (.A(n_1880), .B(n_302), .ZN(n_1881));
   INV_X1 i_1695 (.A(n_1881), .ZN(n_1882));
   OR3_X1 i_1696 (.A1(n_1884), .A2(n_1885), .A3(n_1886), .ZN(n_1883));
   NOR2_X1 i_1697 (.A1(n_325), .A2(n_348), .ZN(n_1884));
   NOR2_X1 i_1698 (.A1(n_302), .A2(n_348), .ZN(n_1885));
   NOR2_X1 i_1699 (.A1(n_302), .A2(n_325), .ZN(n_1886));
   XNOR2_X1 i_1700 (.A(n_279), .B(n_256), .ZN(n_1887));
   XNOR2_X1 i_1701 (.A(n_1887), .B(n_233), .ZN(n_1888));
   INV_X1 i_1702 (.A(n_1888), .ZN(n_1889));
   OR3_X1 i_1703 (.A1(n_1891), .A2(n_1892), .A3(n_1893), .ZN(n_1890));
   NOR2_X1 i_1704 (.A1(n_256), .A2(n_279), .ZN(n_1891));
   NOR2_X1 i_1705 (.A1(n_233), .A2(n_279), .ZN(n_1892));
   NOR2_X1 i_1706 (.A1(n_233), .A2(n_256), .ZN(n_1893));
   XNOR2_X1 i_1707 (.A(n_210), .B(n_187), .ZN(n_1894));
   XNOR2_X1 i_1708 (.A(n_1894), .B(n_164), .ZN(n_1895));
   INV_X1 i_1709 (.A(n_1895), .ZN(n_1896));
   OR3_X1 i_1710 (.A1(n_1898), .A2(n_1899), .A3(n_1900), .ZN(n_1897));
   NOR2_X1 i_1711 (.A1(n_187), .A2(n_210), .ZN(n_1898));
   NOR2_X1 i_1712 (.A1(n_164), .A2(n_210), .ZN(n_1899));
   NOR2_X1 i_1713 (.A1(n_164), .A2(n_187), .ZN(n_1900));
   XNOR2_X1 i_1714 (.A(n_141), .B(n_118), .ZN(n_1901));
   XNOR2_X1 i_1715 (.A(n_1901), .B(n_1829), .ZN(n_1902));
   NAND3_X1 i_1716 (.A1(n_1904), .A2(n_1905), .A3(n_1907), .ZN(n_1903));
   OR2_X1 i_1717 (.A1(n_118), .A2(n_141), .ZN(n_1904));
   NAND2_X1 i_1718 (.A1(n_1829), .A2(n_1906), .ZN(n_1905));
   INV_X1 i_1719 (.A(n_141), .ZN(n_1906));
   NAND2_X1 i_1720 (.A1(n_1829), .A2(n_1908), .ZN(n_1907));
   INV_X1 i_1721 (.A(n_118), .ZN(n_1908));
   FA_X1 i_1722 (.A(n_1822), .B(n_1815), .CI(n_1808), .CO(n_1910), .S(n_1909));
   FA_X1 i_1723 (.A(n_1801), .B(n_1794), .CI(n_1787), .CO(n_1912), .S(n_1911));
   FA_X1 i_1724 (.A(n_1836), .B(n_1834), .CI(n_1902), .CO(n_1914), .S(n_1913));
   FA_X1 i_1725 (.A(n_1896), .B(n_1889), .CI(n_1882), .CO(n_1916), .S(n_1915));
   FA_X1 i_1726 (.A(n_1875), .B(n_1868), .CI(n_1861), .CO(n_1918), .S(n_1917));
   FA_X1 i_1727 (.A(n_1838), .B(n_1911), .CI(n_1909), .CO(n_1920), .S(n_1919));
   FA_X1 i_1728 (.A(n_1842), .B(n_1840), .CI(n_1913), .CO(n_1922), .S(n_1921));
   FA_X1 i_1729 (.A(n_1846), .B(n_1844), .CI(n_1917), .CO(n_1924), .S(n_1923));
   FA_X1 i_1730 (.A(n_1915), .B(n_1848), .CI(n_1921), .CO(n_1926), .S(n_1925));
   FA_X1 i_1731 (.A(n_1919), .B(n_1850), .CI(n_1923), .CO(n_1928), .S(n_1927));
   FA_X1 i_1732 (.A(n_1852), .B(n_1925), .CI(n_1854), .CO(n_1930), .S(n_1929));
   FA_X1 i_1733 (.A(n_1927), .B(n_1856), .CI(n_1929), .CO(n_1932), .S(n_1931));
   XNOR2_X1 i_1734 (.A(n_556), .B(n_533), .ZN(n_1933));
   XNOR2_X1 i_1735 (.A(n_1933), .B(n_510), .ZN(n_1934));
   INV_X1 i_1736 (.A(n_1934), .ZN(n_1935));
   OR3_X1 i_1737 (.A1(n_1937), .A2(n_1938), .A3(n_1939), .ZN(n_1936));
   NOR2_X1 i_1738 (.A1(n_533), .A2(n_556), .ZN(n_1937));
   NOR2_X1 i_1739 (.A1(n_510), .A2(n_556), .ZN(n_1938));
   NOR2_X1 i_1740 (.A1(n_510), .A2(n_533), .ZN(n_1939));
   XNOR2_X1 i_1741 (.A(n_487), .B(n_464), .ZN(n_1940));
   XNOR2_X1 i_1742 (.A(n_1940), .B(n_441), .ZN(n_1941));
   INV_X1 i_1743 (.A(n_1941), .ZN(n_1942));
   OR3_X1 i_1744 (.A1(n_1944), .A2(n_1945), .A3(n_1946), .ZN(n_1943));
   NOR2_X1 i_1745 (.A1(n_464), .A2(n_487), .ZN(n_1944));
   NOR2_X1 i_1746 (.A1(n_441), .A2(n_487), .ZN(n_1945));
   NOR2_X1 i_1747 (.A1(n_441), .A2(n_464), .ZN(n_1946));
   XNOR2_X1 i_1748 (.A(n_418), .B(n_395), .ZN(n_1947));
   XNOR2_X1 i_1749 (.A(n_1947), .B(n_372), .ZN(n_1948));
   INV_X1 i_1750 (.A(n_1948), .ZN(n_1949));
   OR3_X1 i_1751 (.A1(n_1951), .A2(n_1952), .A3(n_1953), .ZN(n_1950));
   NOR2_X1 i_1752 (.A1(n_395), .A2(n_418), .ZN(n_1951));
   NOR2_X1 i_1753 (.A1(n_372), .A2(n_418), .ZN(n_1952));
   NOR2_X1 i_1754 (.A1(n_372), .A2(n_395), .ZN(n_1953));
   XNOR2_X1 i_1755 (.A(n_349), .B(n_326), .ZN(n_1954));
   XNOR2_X1 i_1756 (.A(n_1954), .B(n_303), .ZN(n_1955));
   INV_X1 i_1757 (.A(n_1955), .ZN(n_1956));
   OR3_X1 i_1758 (.A1(n_1958), .A2(n_1959), .A3(n_1960), .ZN(n_1957));
   NOR2_X1 i_1759 (.A1(n_326), .A2(n_349), .ZN(n_1958));
   NOR2_X1 i_1760 (.A1(n_303), .A2(n_349), .ZN(n_1959));
   NOR2_X1 i_1761 (.A1(n_303), .A2(n_326), .ZN(n_1960));
   XNOR2_X1 i_1762 (.A(n_280), .B(n_257), .ZN(n_1961));
   XNOR2_X1 i_1763 (.A(n_1961), .B(n_234), .ZN(n_1962));
   INV_X1 i_1764 (.A(n_1962), .ZN(n_1963));
   OR3_X1 i_1765 (.A1(n_1965), .A2(n_1966), .A3(n_1967), .ZN(n_1964));
   NOR2_X1 i_1766 (.A1(n_257), .A2(n_280), .ZN(n_1965));
   NOR2_X1 i_1767 (.A1(n_234), .A2(n_280), .ZN(n_1966));
   NOR2_X1 i_1768 (.A1(n_234), .A2(n_257), .ZN(n_1967));
   XNOR2_X1 i_1769 (.A(n_211), .B(n_188), .ZN(n_1968));
   XNOR2_X1 i_1770 (.A(n_1968), .B(n_165), .ZN(n_1969));
   INV_X1 i_1771 (.A(n_1969), .ZN(n_1970));
   OR3_X1 i_1772 (.A1(n_1972), .A2(n_1973), .A3(n_1974), .ZN(n_1971));
   NOR2_X1 i_1773 (.A1(n_188), .A2(n_211), .ZN(n_1972));
   NOR2_X1 i_1774 (.A1(n_165), .A2(n_211), .ZN(n_1973));
   NOR2_X1 i_1775 (.A1(n_165), .A2(n_188), .ZN(n_1974));
   XNOR2_X1 i_1776 (.A(n_142), .B(n_1897), .ZN(n_1975));
   XNOR2_X1 i_1777 (.A(n_1975), .B(n_1890), .ZN(n_1976));
   INV_X1 i_1778 (.A(n_1976), .ZN(n_1977));
   NAND3_X1 i_1779 (.A1(n_1979), .A2(n_1981), .A3(n_1982), .ZN(n_1978));
   NAND2_X1 i_1780 (.A1(n_1897), .A2(n_1980), .ZN(n_1979));
   INV_X1 i_1781 (.A(n_142), .ZN(n_1980));
   NAND2_X1 i_1782 (.A1(n_1890), .A2(n_1980), .ZN(n_1981));
   NAND2_X1 i_1783 (.A1(n_1890), .A2(n_1897), .ZN(n_1982));
   FA_X1 i_1784 (.A(n_1883), .B(n_1876), .CI(n_1869), .CO(n_1984), .S(n_1983));
   FA_X1 i_1785 (.A(n_1862), .B(n_1912), .CI(n_1910), .CO(n_1986), .S(n_1985));
   FA_X1 i_1786 (.A(n_1903), .B(n_1970), .CI(n_1963), .CO(n_1988), .S(n_1987));
   FA_X1 i_1787 (.A(n_1956), .B(n_1949), .CI(n_1942), .CO(n_1990), .S(n_1989));
   FA_X1 i_1788 (.A(n_1935), .B(n_1983), .CI(n_1977), .CO(n_1992), .S(n_1991));
   FA_X1 i_1789 (.A(n_1918), .B(n_1916), .CI(n_1914), .CO(n_1994), .S(n_1993));
   FA_X1 i_1790 (.A(n_1985), .B(n_1920), .CI(n_1989), .CO(n_1996), .S(n_1995));
   FA_X1 i_1791 (.A(n_1987), .B(n_1922), .CI(n_1993), .CO(n_1998), .S(n_1997));
   FA_X1 i_1792 (.A(n_1991), .B(n_1924), .CI(n_1995), .CO(n_2000), .S(n_1999));
   FA_X1 i_1793 (.A(n_1926), .B(n_1997), .CI(n_1928), .CO(n_2002), .S(n_2001));
   FA_X1 i_1794 (.A(n_1999), .B(n_1930), .CI(n_2001), .CO(n_2004), .S(n_2003));
   XNOR2_X1 i_1795 (.A(n_557), .B(n_534), .ZN(n_2005));
   XNOR2_X1 i_1796 (.A(n_2005), .B(n_511), .ZN(n_2006));
   INV_X1 i_1797 (.A(n_2006), .ZN(n_2007));
   OR3_X1 i_1798 (.A1(n_2009), .A2(n_2010), .A3(n_2011), .ZN(n_2008));
   NOR2_X1 i_1799 (.A1(n_534), .A2(n_557), .ZN(n_2009));
   NOR2_X1 i_1800 (.A1(n_511), .A2(n_557), .ZN(n_2010));
   NOR2_X1 i_1801 (.A1(n_511), .A2(n_534), .ZN(n_2011));
   XNOR2_X1 i_1802 (.A(n_488), .B(n_465), .ZN(n_2012));
   XNOR2_X1 i_1803 (.A(n_2012), .B(n_442), .ZN(n_2013));
   INV_X1 i_1804 (.A(n_2013), .ZN(n_2014));
   OR3_X1 i_1805 (.A1(n_2016), .A2(n_2017), .A3(n_2018), .ZN(n_2015));
   NOR2_X1 i_1806 (.A1(n_465), .A2(n_488), .ZN(n_2016));
   NOR2_X1 i_1807 (.A1(n_442), .A2(n_488), .ZN(n_2017));
   NOR2_X1 i_1808 (.A1(n_442), .A2(n_465), .ZN(n_2018));
   XNOR2_X1 i_1809 (.A(n_419), .B(n_396), .ZN(n_2019));
   XNOR2_X1 i_1810 (.A(n_2019), .B(n_373), .ZN(n_2020));
   INV_X1 i_1811 (.A(n_2020), .ZN(n_2021));
   OR3_X1 i_1812 (.A1(n_2023), .A2(n_2024), .A3(n_2025), .ZN(n_2022));
   NOR2_X1 i_1813 (.A1(n_396), .A2(n_419), .ZN(n_2023));
   NOR2_X1 i_1814 (.A1(n_373), .A2(n_419), .ZN(n_2024));
   NOR2_X1 i_1815 (.A1(n_373), .A2(n_396), .ZN(n_2025));
   XNOR2_X1 i_1816 (.A(n_350), .B(n_327), .ZN(n_2026));
   XNOR2_X1 i_1817 (.A(n_2026), .B(n_304), .ZN(n_2027));
   INV_X1 i_1818 (.A(n_2027), .ZN(n_2028));
   OR3_X1 i_1819 (.A1(n_2030), .A2(n_2031), .A3(n_2032), .ZN(n_2029));
   NOR2_X1 i_1820 (.A1(n_327), .A2(n_350), .ZN(n_2030));
   NOR2_X1 i_1821 (.A1(n_304), .A2(n_350), .ZN(n_2031));
   NOR2_X1 i_1822 (.A1(n_304), .A2(n_327), .ZN(n_2032));
   XNOR2_X1 i_1823 (.A(n_281), .B(n_258), .ZN(n_2033));
   XNOR2_X1 i_1824 (.A(n_2033), .B(n_235), .ZN(n_2034));
   INV_X1 i_1825 (.A(n_2034), .ZN(n_2035));
   OR3_X1 i_1826 (.A1(n_2037), .A2(n_2038), .A3(n_2039), .ZN(n_2036));
   NOR2_X1 i_1827 (.A1(n_258), .A2(n_281), .ZN(n_2037));
   NOR2_X1 i_1828 (.A1(n_235), .A2(n_281), .ZN(n_2038));
   NOR2_X1 i_1829 (.A1(n_235), .A2(n_258), .ZN(n_2039));
   XNOR2_X1 i_1830 (.A(n_212), .B(n_189), .ZN(n_2040));
   XNOR2_X1 i_1831 (.A(n_2040), .B(n_166), .ZN(n_2041));
   INV_X1 i_1832 (.A(n_2041), .ZN(n_2042));
   OR3_X1 i_1833 (.A1(n_2044), .A2(n_2045), .A3(n_2046), .ZN(n_2043));
   NOR2_X1 i_1834 (.A1(n_189), .A2(n_212), .ZN(n_2044));
   NOR2_X1 i_1835 (.A1(n_166), .A2(n_212), .ZN(n_2045));
   NOR2_X1 i_1836 (.A1(n_166), .A2(n_189), .ZN(n_2046));
   FA_X1 i_1837 (.A(n_1971), .B(n_1964), .CI(n_1957), .CO(n_2048), .S(n_2047));
   FA_X1 i_1838 (.A(n_1950), .B(n_1943), .CI(n_1936), .CO(n_2050), .S(n_2049));
   FA_X1 i_1839 (.A(n_1984), .B(n_1978), .CI(n_2042), .CO(n_2052), .S(n_2051));
   FA_X1 i_1840 (.A(n_2035), .B(n_2028), .CI(n_2021), .CO(n_2054), .S(n_2053));
   FA_X1 i_1841 (.A(n_2014), .B(n_2007), .CI(n_1986), .CO(n_2056), .S(n_2055));
   FA_X1 i_1842 (.A(n_2049), .B(n_2047), .CI(n_1990), .CO(n_2058), .S(n_2057));
   FA_X1 i_1843 (.A(n_1988), .B(n_2051), .CI(n_1994), .CO(n_2060), .S(n_2059));
   FA_X1 i_1844 (.A(n_1992), .B(n_2055), .CI(n_2053), .CO(n_2062), .S(n_2061));
   FA_X1 i_1845 (.A(n_2057), .B(n_1996), .CI(n_2059), .CO(n_2064), .S(n_2063));
   FA_X1 i_1846 (.A(n_1998), .B(n_2061), .CI(n_2000), .CO(n_2066), .S(n_2065));
   FA_X1 i_1847 (.A(n_2063), .B(n_2002), .CI(n_2065), .CO(n_2068), .S(n_2067));
   XNOR2_X1 i_1848 (.A(n_558), .B(n_535), .ZN(n_2069));
   XNOR2_X1 i_1849 (.A(n_2069), .B(n_512), .ZN(n_2070));
   INV_X1 i_1850 (.A(n_2070), .ZN(n_2071));
   OR3_X1 i_1851 (.A1(n_2073), .A2(n_2074), .A3(n_2075), .ZN(n_2072));
   NOR2_X1 i_1852 (.A1(n_535), .A2(n_558), .ZN(n_2073));
   NOR2_X1 i_1853 (.A1(n_512), .A2(n_558), .ZN(n_2074));
   NOR2_X1 i_1854 (.A1(n_512), .A2(n_535), .ZN(n_2075));
   XNOR2_X1 i_1855 (.A(n_489), .B(n_466), .ZN(n_2076));
   XNOR2_X1 i_1856 (.A(n_2076), .B(n_443), .ZN(n_2077));
   INV_X1 i_1857 (.A(n_2077), .ZN(n_2078));
   OR3_X1 i_1858 (.A1(n_2080), .A2(n_2081), .A3(n_2082), .ZN(n_2079));
   NOR2_X1 i_1859 (.A1(n_466), .A2(n_489), .ZN(n_2080));
   NOR2_X1 i_1860 (.A1(n_443), .A2(n_489), .ZN(n_2081));
   NOR2_X1 i_1861 (.A1(n_443), .A2(n_466), .ZN(n_2082));
   XNOR2_X1 i_1862 (.A(n_420), .B(n_397), .ZN(n_2083));
   XNOR2_X1 i_1863 (.A(n_2083), .B(n_374), .ZN(n_2084));
   INV_X1 i_1864 (.A(n_2084), .ZN(n_2085));
   OR3_X1 i_1865 (.A1(n_2087), .A2(n_2088), .A3(n_2089), .ZN(n_2086));
   NOR2_X1 i_1866 (.A1(n_397), .A2(n_420), .ZN(n_2087));
   NOR2_X1 i_1867 (.A1(n_374), .A2(n_420), .ZN(n_2088));
   NOR2_X1 i_1868 (.A1(n_374), .A2(n_397), .ZN(n_2089));
   XNOR2_X1 i_1869 (.A(n_351), .B(n_328), .ZN(n_2090));
   XNOR2_X1 i_1870 (.A(n_2090), .B(n_305), .ZN(n_2091));
   INV_X1 i_1871 (.A(n_2091), .ZN(n_2092));
   OR3_X1 i_1872 (.A1(n_2094), .A2(n_2095), .A3(n_2096), .ZN(n_2093));
   NOR2_X1 i_1873 (.A1(n_328), .A2(n_351), .ZN(n_2094));
   NOR2_X1 i_1874 (.A1(n_305), .A2(n_351), .ZN(n_2095));
   NOR2_X1 i_1875 (.A1(n_305), .A2(n_328), .ZN(n_2096));
   XNOR2_X1 i_1876 (.A(n_282), .B(n_259), .ZN(n_2097));
   XNOR2_X1 i_1877 (.A(n_2097), .B(n_236), .ZN(n_2098));
   INV_X1 i_1878 (.A(n_2098), .ZN(n_2099));
   OR3_X1 i_1879 (.A1(n_2101), .A2(n_2102), .A3(n_2103), .ZN(n_2100));
   NOR2_X1 i_1880 (.A1(n_259), .A2(n_282), .ZN(n_2101));
   NOR2_X1 i_1881 (.A1(n_236), .A2(n_282), .ZN(n_2102));
   NOR2_X1 i_1882 (.A1(n_236), .A2(n_259), .ZN(n_2103));
   XNOR2_X1 i_1883 (.A(n_213), .B(n_190), .ZN(n_2104));
   XNOR2_X1 i_1884 (.A(n_2104), .B(n_2043), .ZN(n_2105));
   NAND3_X1 i_1885 (.A1(n_2107), .A2(n_2108), .A3(n_2110), .ZN(n_2106));
   OR2_X1 i_1886 (.A1(n_190), .A2(n_213), .ZN(n_2107));
   NAND2_X1 i_1887 (.A1(n_2043), .A2(n_2109), .ZN(n_2108));
   INV_X1 i_1888 (.A(n_213), .ZN(n_2109));
   NAND2_X1 i_1889 (.A1(n_2043), .A2(n_2111), .ZN(n_2110));
   INV_X1 i_1890 (.A(n_190), .ZN(n_2111));
   FA_X1 i_1891 (.A(n_2036), .B(n_2029), .CI(n_2022), .CO(n_2113), .S(n_2112));
   FA_X1 i_1892 (.A(n_2015), .B(n_2008), .CI(n_2050), .CO(n_2115), .S(n_2114));
   FA_X1 i_1893 (.A(n_2048), .B(n_2105), .CI(n_2099), .CO(n_2117), .S(n_2116));
   FA_X1 i_1894 (.A(n_2092), .B(n_2085), .CI(n_2078), .CO(n_2119), .S(n_2118));
   FA_X1 i_1895 (.A(n_2071), .B(n_2114), .CI(n_2112), .CO(n_2121), .S(n_2120));
   FA_X1 i_1896 (.A(n_2054), .B(n_2052), .CI(n_2056), .CO(n_2123), .S(n_2122));
   FA_X1 i_1897 (.A(n_2058), .B(n_2118), .CI(n_2116), .CO(n_2125), .S(n_2124));
   FA_X1 i_1898 (.A(n_2060), .B(n_2122), .CI(n_2120), .CO(n_2127), .S(n_2126));
   FA_X1 i_1899 (.A(n_2062), .B(n_2124), .CI(n_2064), .CO(n_2129), .S(n_2128));
   FA_X1 i_1900 (.A(n_2126), .B(n_2066), .CI(n_2128), .CO(n_2131), .S(n_2130));
   XNOR2_X1 i_1901 (.A(n_559), .B(n_536), .ZN(n_2132));
   XNOR2_X1 i_1902 (.A(n_2132), .B(n_513), .ZN(n_2133));
   INV_X1 i_1903 (.A(n_2133), .ZN(n_2134));
   OR3_X1 i_1904 (.A1(n_2136), .A2(n_2137), .A3(n_2138), .ZN(n_2135));
   NOR2_X1 i_1905 (.A1(n_536), .A2(n_559), .ZN(n_2136));
   NOR2_X1 i_1906 (.A1(n_513), .A2(n_559), .ZN(n_2137));
   NOR2_X1 i_1907 (.A1(n_513), .A2(n_536), .ZN(n_2138));
   XNOR2_X1 i_1908 (.A(n_490), .B(n_467), .ZN(n_2139));
   XNOR2_X1 i_1909 (.A(n_2139), .B(n_444), .ZN(n_2140));
   INV_X1 i_1910 (.A(n_2140), .ZN(n_2141));
   OR3_X1 i_1911 (.A1(n_2143), .A2(n_2144), .A3(n_2145), .ZN(n_2142));
   NOR2_X1 i_1912 (.A1(n_467), .A2(n_490), .ZN(n_2143));
   NOR2_X1 i_1913 (.A1(n_444), .A2(n_490), .ZN(n_2144));
   NOR2_X1 i_1914 (.A1(n_444), .A2(n_467), .ZN(n_2145));
   XNOR2_X1 i_1915 (.A(n_421), .B(n_398), .ZN(n_2146));
   XNOR2_X1 i_1916 (.A(n_2146), .B(n_375), .ZN(n_2147));
   INV_X1 i_1917 (.A(n_2147), .ZN(n_2148));
   OR3_X1 i_1918 (.A1(n_2150), .A2(n_2151), .A3(n_2152), .ZN(n_2149));
   NOR2_X1 i_1919 (.A1(n_398), .A2(n_421), .ZN(n_2150));
   NOR2_X1 i_1920 (.A1(n_375), .A2(n_421), .ZN(n_2151));
   NOR2_X1 i_1921 (.A1(n_375), .A2(n_398), .ZN(n_2152));
   XNOR2_X1 i_1922 (.A(n_352), .B(n_329), .ZN(n_2153));
   XNOR2_X1 i_1923 (.A(n_2153), .B(n_306), .ZN(n_2154));
   INV_X1 i_1924 (.A(n_2154), .ZN(n_2155));
   OR3_X1 i_1925 (.A1(n_2157), .A2(n_2158), .A3(n_2159), .ZN(n_2156));
   NOR2_X1 i_1926 (.A1(n_329), .A2(n_352), .ZN(n_2157));
   NOR2_X1 i_1927 (.A1(n_306), .A2(n_352), .ZN(n_2158));
   NOR2_X1 i_1928 (.A1(n_306), .A2(n_329), .ZN(n_2159));
   XNOR2_X1 i_1929 (.A(n_283), .B(n_260), .ZN(n_2160));
   XNOR2_X1 i_1930 (.A(n_2160), .B(n_237), .ZN(n_2161));
   INV_X1 i_1931 (.A(n_2161), .ZN(n_2162));
   OR3_X1 i_1932 (.A1(n_2164), .A2(n_2165), .A3(n_2166), .ZN(n_2163));
   NOR2_X1 i_1933 (.A1(n_260), .A2(n_283), .ZN(n_2164));
   NOR2_X1 i_1934 (.A1(n_237), .A2(n_283), .ZN(n_2165));
   NOR2_X1 i_1935 (.A1(n_237), .A2(n_260), .ZN(n_2166));
   XNOR2_X1 i_1936 (.A(n_214), .B(n_2100), .ZN(n_2167));
   XNOR2_X1 i_1937 (.A(n_2167), .B(n_2093), .ZN(n_2168));
   INV_X1 i_1938 (.A(n_2168), .ZN(n_2169));
   NAND3_X1 i_1939 (.A1(n_2171), .A2(n_2173), .A3(n_2174), .ZN(n_2170));
   NAND2_X1 i_1940 (.A1(n_2100), .A2(n_2172), .ZN(n_2171));
   INV_X1 i_1941 (.A(n_214), .ZN(n_2172));
   NAND2_X1 i_1942 (.A1(n_2093), .A2(n_2172), .ZN(n_2173));
   NAND2_X1 i_1943 (.A1(n_2093), .A2(n_2100), .ZN(n_2174));
   FA_X1 i_1944 (.A(n_2086), .B(n_2079), .CI(n_2072), .CO(n_2176), .S(n_2175));
   FA_X1 i_1945 (.A(n_2113), .B(n_2106), .CI(n_2162), .CO(n_2178), .S(n_2177));
   FA_X1 i_1946 (.A(n_2155), .B(n_2148), .CI(n_2141), .CO(n_2180), .S(n_2179));
   FA_X1 i_1947 (.A(n_2134), .B(n_2115), .CI(n_2175), .CO(n_2182), .S(n_2181));
   FA_X1 i_1948 (.A(n_2169), .B(n_2119), .CI(n_2117), .CO(n_2184), .S(n_2183));
   FA_X1 i_1949 (.A(n_2177), .B(n_2121), .CI(n_2123), .CO(n_2186), .S(n_2185));
   FA_X1 i_1950 (.A(n_2179), .B(n_2181), .CI(n_2183), .CO(n_2188), .S(n_2187));
   FA_X1 i_1951 (.A(n_2125), .B(n_2185), .CI(n_2127), .CO(n_2190), .S(n_2189));
   FA_X1 i_1952 (.A(n_2187), .B(n_2129), .CI(n_2189), .CO(n_2192), .S(n_2191));
   XNOR2_X1 i_1953 (.A(n_560), .B(n_537), .ZN(n_2193));
   XNOR2_X1 i_1954 (.A(n_2193), .B(n_514), .ZN(n_2194));
   INV_X1 i_1955 (.A(n_2194), .ZN(n_2195));
   OR3_X1 i_1956 (.A1(n_2197), .A2(n_2198), .A3(n_2199), .ZN(n_2196));
   NOR2_X1 i_1957 (.A1(n_537), .A2(n_560), .ZN(n_2197));
   NOR2_X1 i_1958 (.A1(n_514), .A2(n_560), .ZN(n_2198));
   NOR2_X1 i_1959 (.A1(n_514), .A2(n_537), .ZN(n_2199));
   XNOR2_X1 i_1960 (.A(n_491), .B(n_468), .ZN(n_2200));
   XNOR2_X1 i_1961 (.A(n_2200), .B(n_445), .ZN(n_2201));
   INV_X1 i_1962 (.A(n_2201), .ZN(n_2202));
   OR3_X1 i_1963 (.A1(n_2204), .A2(n_2205), .A3(n_2206), .ZN(n_2203));
   NOR2_X1 i_1964 (.A1(n_468), .A2(n_491), .ZN(n_2204));
   NOR2_X1 i_1965 (.A1(n_445), .A2(n_491), .ZN(n_2205));
   NOR2_X1 i_1966 (.A1(n_445), .A2(n_468), .ZN(n_2206));
   XNOR2_X1 i_1967 (.A(n_422), .B(n_399), .ZN(n_2207));
   XNOR2_X1 i_1968 (.A(n_2207), .B(n_376), .ZN(n_2208));
   INV_X1 i_1969 (.A(n_2208), .ZN(n_2209));
   OR3_X1 i_1970 (.A1(n_2211), .A2(n_2212), .A3(n_2213), .ZN(n_2210));
   NOR2_X1 i_1971 (.A1(n_399), .A2(n_422), .ZN(n_2211));
   NOR2_X1 i_1972 (.A1(n_376), .A2(n_422), .ZN(n_2212));
   NOR2_X1 i_1973 (.A1(n_376), .A2(n_399), .ZN(n_2213));
   XNOR2_X1 i_1974 (.A(n_353), .B(n_330), .ZN(n_2214));
   XNOR2_X1 i_1975 (.A(n_2214), .B(n_307), .ZN(n_2215));
   INV_X1 i_1976 (.A(n_2215), .ZN(n_2216));
   OR3_X1 i_1977 (.A1(n_2218), .A2(n_2219), .A3(n_2220), .ZN(n_2217));
   NOR2_X1 i_1978 (.A1(n_330), .A2(n_353), .ZN(n_2218));
   NOR2_X1 i_1979 (.A1(n_307), .A2(n_353), .ZN(n_2219));
   NOR2_X1 i_1980 (.A1(n_307), .A2(n_330), .ZN(n_2220));
   XNOR2_X1 i_1981 (.A(n_284), .B(n_261), .ZN(n_2221));
   XNOR2_X1 i_1982 (.A(n_2221), .B(n_238), .ZN(n_2222));
   INV_X1 i_1983 (.A(n_2222), .ZN(n_2223));
   OR3_X1 i_1984 (.A1(n_2225), .A2(n_2226), .A3(n_2227), .ZN(n_2224));
   NOR2_X1 i_1985 (.A1(n_261), .A2(n_284), .ZN(n_2225));
   NOR2_X1 i_1986 (.A1(n_238), .A2(n_284), .ZN(n_2226));
   NOR2_X1 i_1987 (.A1(n_238), .A2(n_261), .ZN(n_2227));
   FA_X1 i_1988 (.A(n_2163), .B(n_2156), .CI(n_2149), .CO(n_2229), .S(n_2228));
   FA_X1 i_1989 (.A(n_2142), .B(n_2135), .CI(n_2176), .CO(n_2231), .S(n_2230));
   FA_X1 i_1990 (.A(n_2170), .B(n_2223), .CI(n_2216), .CO(n_2233), .S(n_2232));
   FA_X1 i_1991 (.A(n_2209), .B(n_2202), .CI(n_2195), .CO(n_2235), .S(n_2234));
   FA_X1 i_1992 (.A(n_2230), .B(n_2228), .CI(n_2180), .CO(n_2237), .S(n_2236));
   FA_X1 i_1993 (.A(n_2178), .B(n_2184), .CI(n_2182), .CO(n_2239), .S(n_2238));
   FA_X1 i_1994 (.A(n_2234), .B(n_2232), .CI(n_2186), .CO(n_2241), .S(n_2240));
   FA_X1 i_1995 (.A(n_2236), .B(n_2238), .CI(n_2188), .CO(n_2243), .S(n_2242));
   FA_X1 i_1996 (.A(n_2240), .B(n_2190), .CI(n_2242), .CO(n_2245), .S(n_2244));
   XNOR2_X1 i_1997 (.A(n_561), .B(n_538), .ZN(n_2246));
   XNOR2_X1 i_1998 (.A(n_2246), .B(n_515), .ZN(n_2247));
   INV_X1 i_1999 (.A(n_2247), .ZN(n_2248));
   OR3_X1 i_2000 (.A1(n_2250), .A2(n_2251), .A3(n_2252), .ZN(n_2249));
   NOR2_X1 i_2001 (.A1(n_538), .A2(n_561), .ZN(n_2250));
   NOR2_X1 i_2002 (.A1(n_515), .A2(n_561), .ZN(n_2251));
   NOR2_X1 i_2003 (.A1(n_515), .A2(n_538), .ZN(n_2252));
   XNOR2_X1 i_2004 (.A(n_492), .B(n_469), .ZN(n_2253));
   XNOR2_X1 i_2005 (.A(n_2253), .B(n_446), .ZN(n_2254));
   INV_X1 i_2006 (.A(n_2254), .ZN(n_2255));
   OR3_X1 i_2007 (.A1(n_2257), .A2(n_2258), .A3(n_2259), .ZN(n_2256));
   NOR2_X1 i_2008 (.A1(n_469), .A2(n_492), .ZN(n_2257));
   NOR2_X1 i_2009 (.A1(n_446), .A2(n_492), .ZN(n_2258));
   NOR2_X1 i_2010 (.A1(n_446), .A2(n_469), .ZN(n_2259));
   XNOR2_X1 i_2011 (.A(n_423), .B(n_400), .ZN(n_2260));
   XNOR2_X1 i_2012 (.A(n_2260), .B(n_377), .ZN(n_2261));
   INV_X1 i_2013 (.A(n_2261), .ZN(n_2262));
   OR3_X1 i_2014 (.A1(n_2264), .A2(n_2265), .A3(n_2266), .ZN(n_2263));
   NOR2_X1 i_2015 (.A1(n_400), .A2(n_423), .ZN(n_2264));
   NOR2_X1 i_2016 (.A1(n_377), .A2(n_423), .ZN(n_2265));
   NOR2_X1 i_2017 (.A1(n_377), .A2(n_400), .ZN(n_2266));
   XNOR2_X1 i_2018 (.A(n_354), .B(n_331), .ZN(n_2267));
   XNOR2_X1 i_2019 (.A(n_2267), .B(n_308), .ZN(n_2268));
   INV_X1 i_2020 (.A(n_2268), .ZN(n_2269));
   OR3_X1 i_2021 (.A1(n_2271), .A2(n_2272), .A3(n_2273), .ZN(n_2270));
   NOR2_X1 i_2022 (.A1(n_331), .A2(n_354), .ZN(n_2271));
   NOR2_X1 i_2023 (.A1(n_308), .A2(n_354), .ZN(n_2272));
   NOR2_X1 i_2024 (.A1(n_308), .A2(n_331), .ZN(n_2273));
   XNOR2_X1 i_2025 (.A(n_285), .B(n_262), .ZN(n_2274));
   XNOR2_X1 i_2026 (.A(n_2274), .B(n_2224), .ZN(n_2275));
   NAND3_X1 i_2027 (.A1(n_2277), .A2(n_2278), .A3(n_2280), .ZN(n_2276));
   OR2_X1 i_2028 (.A1(n_262), .A2(n_285), .ZN(n_2277));
   NAND2_X1 i_2029 (.A1(n_2224), .A2(n_2279), .ZN(n_2278));
   INV_X1 i_2030 (.A(n_285), .ZN(n_2279));
   NAND2_X1 i_2031 (.A1(n_2224), .A2(n_2281), .ZN(n_2280));
   INV_X1 i_2032 (.A(n_262), .ZN(n_2281));
   FA_X1 i_2033 (.A(n_2217), .B(n_2210), .CI(n_2203), .CO(n_2283), .S(n_2282));
   FA_X1 i_2034 (.A(n_2196), .B(n_2229), .CI(n_2275), .CO(n_2285), .S(n_2284));
   FA_X1 i_2035 (.A(n_2269), .B(n_2262), .CI(n_2255), .CO(n_2287), .S(n_2286));
   FA_X1 i_2036 (.A(n_2248), .B(n_2231), .CI(n_2282), .CO(n_2289), .S(n_2288));
   FA_X1 i_2037 (.A(n_2235), .B(n_2233), .CI(n_2284), .CO(n_2291), .S(n_2290));
   FA_X1 i_2038 (.A(n_2237), .B(n_2286), .CI(n_2288), .CO(n_2293), .S(n_2292));
   FA_X1 i_2039 (.A(n_2239), .B(n_2290), .CI(n_2241), .CO(n_2295), .S(n_2294));
   FA_X1 i_2040 (.A(n_2292), .B(n_2243), .CI(n_2294), .CO(n_2297), .S(n_2296));
   XNOR2_X1 i_2041 (.A(n_562), .B(n_539), .ZN(n_2298));
   XNOR2_X1 i_2042 (.A(n_2298), .B(n_516), .ZN(n_2299));
   INV_X1 i_2043 (.A(n_2299), .ZN(n_2300));
   OR3_X1 i_2044 (.A1(n_2302), .A2(n_2303), .A3(n_2304), .ZN(n_2301));
   NOR2_X1 i_2045 (.A1(n_539), .A2(n_562), .ZN(n_2302));
   NOR2_X1 i_2046 (.A1(n_516), .A2(n_562), .ZN(n_2303));
   NOR2_X1 i_2047 (.A1(n_516), .A2(n_539), .ZN(n_2304));
   XNOR2_X1 i_2048 (.A(n_493), .B(n_470), .ZN(n_2305));
   XNOR2_X1 i_2049 (.A(n_2305), .B(n_447), .ZN(n_2306));
   INV_X1 i_2050 (.A(n_2306), .ZN(n_2307));
   OR3_X1 i_2051 (.A1(n_2309), .A2(n_2310), .A3(n_2311), .ZN(n_2308));
   NOR2_X1 i_2052 (.A1(n_470), .A2(n_493), .ZN(n_2309));
   NOR2_X1 i_2053 (.A1(n_447), .A2(n_493), .ZN(n_2310));
   NOR2_X1 i_2054 (.A1(n_447), .A2(n_470), .ZN(n_2311));
   XNOR2_X1 i_2055 (.A(n_424), .B(n_401), .ZN(n_2312));
   XNOR2_X1 i_2056 (.A(n_2312), .B(n_378), .ZN(n_2313));
   INV_X1 i_2057 (.A(n_2313), .ZN(n_2314));
   OR3_X1 i_2058 (.A1(n_2316), .A2(n_2317), .A3(n_2318), .ZN(n_2315));
   NOR2_X1 i_2059 (.A1(n_401), .A2(n_424), .ZN(n_2316));
   NOR2_X1 i_2060 (.A1(n_378), .A2(n_424), .ZN(n_2317));
   NOR2_X1 i_2061 (.A1(n_378), .A2(n_401), .ZN(n_2318));
   XNOR2_X1 i_2062 (.A(n_355), .B(n_332), .ZN(n_2319));
   XNOR2_X1 i_2063 (.A(n_2319), .B(n_309), .ZN(n_2320));
   INV_X1 i_2064 (.A(n_2320), .ZN(n_2321));
   OR3_X1 i_2065 (.A1(n_2323), .A2(n_2324), .A3(n_2325), .ZN(n_2322));
   NOR2_X1 i_2066 (.A1(n_332), .A2(n_355), .ZN(n_2323));
   NOR2_X1 i_2067 (.A1(n_309), .A2(n_355), .ZN(n_2324));
   NOR2_X1 i_2068 (.A1(n_309), .A2(n_332), .ZN(n_2325));
   XNOR2_X1 i_2069 (.A(n_286), .B(n_2270), .ZN(n_2326));
   XNOR2_X1 i_2070 (.A(n_2326), .B(n_2263), .ZN(n_2327));
   INV_X1 i_2071 (.A(n_2327), .ZN(n_2328));
   NAND3_X1 i_2072 (.A1(n_2330), .A2(n_2332), .A3(n_2333), .ZN(n_2329));
   NAND2_X1 i_2073 (.A1(n_2270), .A2(n_2331), .ZN(n_2330));
   INV_X1 i_2074 (.A(n_286), .ZN(n_2331));
   NAND2_X1 i_2075 (.A1(n_2263), .A2(n_2331), .ZN(n_2332));
   NAND2_X1 i_2076 (.A1(n_2263), .A2(n_2270), .ZN(n_2333));
   FA_X1 i_2077 (.A(n_2256), .B(n_2249), .CI(n_2283), .CO(n_2335), .S(n_2334));
   FA_X1 i_2078 (.A(n_2276), .B(n_2321), .CI(n_2314), .CO(n_2337), .S(n_2336));
   FA_X1 i_2079 (.A(n_2307), .B(n_2300), .CI(n_2334), .CO(n_2339), .S(n_2338));
   FA_X1 i_2080 (.A(n_2328), .B(n_2287), .CI(n_2285), .CO(n_2341), .S(n_2340));
   FA_X1 i_2081 (.A(n_2289), .B(n_2338), .CI(n_2336), .CO(n_2343), .S(n_2342));
   FA_X1 i_2082 (.A(n_2291), .B(n_2340), .CI(n_2293), .CO(n_2345), .S(n_2344));
   FA_X1 i_2083 (.A(n_2295), .B(n_2342), .CI(n_2344), .CO(n_2347), .S(n_2346));
   XNOR2_X1 i_2084 (.A(n_563), .B(n_540), .ZN(n_2348));
   XNOR2_X1 i_2085 (.A(n_2348), .B(n_517), .ZN(n_2349));
   INV_X1 i_2086 (.A(n_2349), .ZN(n_2350));
   OR3_X1 i_2087 (.A1(n_2352), .A2(n_2353), .A3(n_2354), .ZN(n_2351));
   NOR2_X1 i_2088 (.A1(n_540), .A2(n_563), .ZN(n_2352));
   NOR2_X1 i_2089 (.A1(n_517), .A2(n_563), .ZN(n_2353));
   NOR2_X1 i_2090 (.A1(n_517), .A2(n_540), .ZN(n_2354));
   XNOR2_X1 i_2091 (.A(n_494), .B(n_471), .ZN(n_2355));
   XNOR2_X1 i_2092 (.A(n_2355), .B(n_448), .ZN(n_2356));
   INV_X1 i_2093 (.A(n_2356), .ZN(n_2357));
   OR3_X1 i_2094 (.A1(n_2359), .A2(n_2360), .A3(n_2361), .ZN(n_2358));
   NOR2_X1 i_2095 (.A1(n_471), .A2(n_494), .ZN(n_2359));
   NOR2_X1 i_2096 (.A1(n_448), .A2(n_494), .ZN(n_2360));
   NOR2_X1 i_2097 (.A1(n_448), .A2(n_471), .ZN(n_2361));
   XNOR2_X1 i_2098 (.A(n_425), .B(n_402), .ZN(n_2362));
   XNOR2_X1 i_2099 (.A(n_2362), .B(n_379), .ZN(n_2363));
   INV_X1 i_2100 (.A(n_2363), .ZN(n_2364));
   OR3_X1 i_2101 (.A1(n_2366), .A2(n_2367), .A3(n_2368), .ZN(n_2365));
   NOR2_X1 i_2102 (.A1(n_402), .A2(n_425), .ZN(n_2366));
   NOR2_X1 i_2103 (.A1(n_379), .A2(n_425), .ZN(n_2367));
   NOR2_X1 i_2104 (.A1(n_379), .A2(n_402), .ZN(n_2368));
   XNOR2_X1 i_2105 (.A(n_356), .B(n_333), .ZN(n_2369));
   XNOR2_X1 i_2106 (.A(n_2369), .B(n_310), .ZN(n_2370));
   INV_X1 i_2107 (.A(n_2370), .ZN(n_2371));
   OR3_X1 i_2108 (.A1(n_2373), .A2(n_2374), .A3(n_2375), .ZN(n_2372));
   NOR2_X1 i_2109 (.A1(n_333), .A2(n_356), .ZN(n_2373));
   NOR2_X1 i_2110 (.A1(n_310), .A2(n_356), .ZN(n_2374));
   NOR2_X1 i_2111 (.A1(n_310), .A2(n_333), .ZN(n_2375));
   FA_X1 i_2112 (.A(n_2322), .B(n_2315), .CI(n_2308), .CO(n_2377), .S(n_2376));
   FA_X1 i_2113 (.A(n_2301), .B(n_2329), .CI(n_2371), .CO(n_2379), .S(n_2378));
   FA_X1 i_2114 (.A(n_2364), .B(n_2357), .CI(n_2350), .CO(n_2381), .S(n_2380));
   FA_X1 i_2115 (.A(n_2335), .B(n_2376), .CI(n_2337), .CO(n_2383), .S(n_2382));
   FA_X1 i_2116 (.A(n_2378), .B(n_2341), .CI(n_2339), .CO(n_2385), .S(n_2384));
   FA_X1 i_2117 (.A(n_2380), .B(n_2382), .CI(n_2343), .CO(n_2387), .S(n_2386));
   FA_X1 i_2118 (.A(n_2384), .B(n_2345), .CI(n_2386), .CO(n_2389), .S(n_2388));
   XNOR2_X1 i_2119 (.A(n_564), .B(n_541), .ZN(n_2390));
   XNOR2_X1 i_2120 (.A(n_2390), .B(n_518), .ZN(n_2391));
   INV_X1 i_2121 (.A(n_2391), .ZN(n_2392));
   OR3_X1 i_2122 (.A1(n_2394), .A2(n_2395), .A3(n_2396), .ZN(n_2393));
   NOR2_X1 i_2123 (.A1(n_541), .A2(n_564), .ZN(n_2394));
   NOR2_X1 i_2124 (.A1(n_518), .A2(n_564), .ZN(n_2395));
   NOR2_X1 i_2125 (.A1(n_518), .A2(n_541), .ZN(n_2396));
   XNOR2_X1 i_2126 (.A(n_495), .B(n_472), .ZN(n_2397));
   XNOR2_X1 i_2127 (.A(n_2397), .B(n_449), .ZN(n_2398));
   INV_X1 i_2128 (.A(n_2398), .ZN(n_2399));
   OR3_X1 i_2129 (.A1(n_2401), .A2(n_2402), .A3(n_2403), .ZN(n_2400));
   NOR2_X1 i_2130 (.A1(n_472), .A2(n_495), .ZN(n_2401));
   NOR2_X1 i_2131 (.A1(n_449), .A2(n_495), .ZN(n_2402));
   NOR2_X1 i_2132 (.A1(n_449), .A2(n_472), .ZN(n_2403));
   XNOR2_X1 i_2133 (.A(n_426), .B(n_403), .ZN(n_2404));
   XNOR2_X1 i_2134 (.A(n_2404), .B(n_380), .ZN(n_2405));
   INV_X1 i_2135 (.A(n_2405), .ZN(n_2406));
   OR3_X1 i_2136 (.A1(n_2408), .A2(n_2409), .A3(n_2410), .ZN(n_2407));
   NOR2_X1 i_2137 (.A1(n_403), .A2(n_426), .ZN(n_2408));
   NOR2_X1 i_2138 (.A1(n_380), .A2(n_426), .ZN(n_2409));
   NOR2_X1 i_2139 (.A1(n_380), .A2(n_403), .ZN(n_2410));
   XNOR2_X1 i_2140 (.A(n_357), .B(n_334), .ZN(n_2411));
   XNOR2_X1 i_2141 (.A(n_2411), .B(n_2372), .ZN(n_2412));
   NAND3_X1 i_2142 (.A1(n_2414), .A2(n_2415), .A3(n_2417), .ZN(n_2413));
   OR2_X1 i_2143 (.A1(n_334), .A2(n_357), .ZN(n_2414));
   NAND2_X1 i_2144 (.A1(n_2372), .A2(n_2416), .ZN(n_2415));
   INV_X1 i_2145 (.A(n_357), .ZN(n_2416));
   NAND2_X1 i_2146 (.A1(n_2372), .A2(n_2418), .ZN(n_2417));
   INV_X1 i_2147 (.A(n_334), .ZN(n_2418));
   FA_X1 i_2148 (.A(n_2365), .B(n_2358), .CI(n_2351), .CO(n_2420), .S(n_2419));
   FA_X1 i_2149 (.A(n_2377), .B(n_2412), .CI(n_2406), .CO(n_2422), .S(n_2421));
   FA_X1 i_2150 (.A(n_2399), .B(n_2392), .CI(n_2419), .CO(n_2424), .S(n_2423));
   FA_X1 i_2151 (.A(n_2381), .B(n_2379), .CI(n_2383), .CO(n_2426), .S(n_2425));
   FA_X1 i_2152 (.A(n_2423), .B(n_2421), .CI(n_2385), .CO(n_2428), .S(n_2427));
   FA_X1 i_2153 (.A(n_2425), .B(n_2387), .CI(n_2427), .CO(n_2430), .S(n_2429));
   XNOR2_X1 i_2154 (.A(n_565), .B(n_542), .ZN(n_2431));
   XNOR2_X1 i_2155 (.A(n_2431), .B(n_519), .ZN(n_2432));
   INV_X1 i_2156 (.A(n_2432), .ZN(n_2433));
   OR3_X1 i_2157 (.A1(n_2435), .A2(n_2436), .A3(n_2437), .ZN(n_2434));
   NOR2_X1 i_2158 (.A1(n_542), .A2(n_565), .ZN(n_2435));
   NOR2_X1 i_2159 (.A1(n_519), .A2(n_565), .ZN(n_2436));
   NOR2_X1 i_2160 (.A1(n_519), .A2(n_542), .ZN(n_2437));
   XNOR2_X1 i_2161 (.A(n_496), .B(n_473), .ZN(n_2438));
   XNOR2_X1 i_2162 (.A(n_2438), .B(n_450), .ZN(n_2439));
   INV_X1 i_2163 (.A(n_2439), .ZN(n_2440));
   OR3_X1 i_2164 (.A1(n_2442), .A2(n_2443), .A3(n_2444), .ZN(n_2441));
   NOR2_X1 i_2165 (.A1(n_473), .A2(n_496), .ZN(n_2442));
   NOR2_X1 i_2166 (.A1(n_450), .A2(n_496), .ZN(n_2443));
   NOR2_X1 i_2167 (.A1(n_450), .A2(n_473), .ZN(n_2444));
   XNOR2_X1 i_2168 (.A(n_427), .B(n_404), .ZN(n_2445));
   XNOR2_X1 i_2169 (.A(n_2445), .B(n_381), .ZN(n_2446));
   INV_X1 i_2170 (.A(n_2446), .ZN(n_2447));
   OR3_X1 i_2171 (.A1(n_2449), .A2(n_2450), .A3(n_2451), .ZN(n_2448));
   NOR2_X1 i_2172 (.A1(n_404), .A2(n_427), .ZN(n_2449));
   NOR2_X1 i_2173 (.A1(n_381), .A2(n_427), .ZN(n_2450));
   NOR2_X1 i_2174 (.A1(n_381), .A2(n_404), .ZN(n_2451));
   XNOR2_X1 i_2175 (.A(n_358), .B(n_2407), .ZN(n_2452));
   XNOR2_X1 i_2176 (.A(n_2452), .B(n_2400), .ZN(n_2453));
   INV_X1 i_2177 (.A(n_2453), .ZN(n_2454));
   NAND3_X1 i_2178 (.A1(n_2456), .A2(n_2458), .A3(n_2459), .ZN(n_2455));
   NAND2_X1 i_2179 (.A1(n_2407), .A2(n_2457), .ZN(n_2456));
   INV_X1 i_2180 (.A(n_358), .ZN(n_2457));
   NAND2_X1 i_2181 (.A1(n_2400), .A2(n_2457), .ZN(n_2458));
   NAND2_X1 i_2182 (.A1(n_2400), .A2(n_2407), .ZN(n_2459));
   FA_X1 i_2183 (.A(n_2393), .B(n_2420), .CI(n_2413), .CO(n_2461), .S(n_2460));
   FA_X1 i_2184 (.A(n_2447), .B(n_2440), .CI(n_2433), .CO(n_2463), .S(n_2462));
   FA_X1 i_2185 (.A(n_2454), .B(n_2422), .CI(n_2460), .CO(n_2465), .S(n_2464));
   FA_X1 i_2186 (.A(n_2424), .B(n_2462), .CI(n_2426), .CO(n_2467), .S(n_2466));
   FA_X1 i_2187 (.A(n_2464), .B(n_2428), .CI(n_2466), .CO(n_2469), .S(n_2468));
   XNOR2_X1 i_2188 (.A(n_566), .B(n_543), .ZN(n_2470));
   XNOR2_X1 i_2189 (.A(n_2470), .B(n_520), .ZN(n_2471));
   INV_X1 i_2190 (.A(n_2471), .ZN(n_2472));
   OR3_X1 i_2191 (.A1(n_2474), .A2(n_2475), .A3(n_2476), .ZN(n_2473));
   NOR2_X1 i_2192 (.A1(n_543), .A2(n_566), .ZN(n_2474));
   NOR2_X1 i_2193 (.A1(n_520), .A2(n_566), .ZN(n_2475));
   NOR2_X1 i_2194 (.A1(n_520), .A2(n_543), .ZN(n_2476));
   XNOR2_X1 i_2195 (.A(n_497), .B(n_474), .ZN(n_2477));
   XNOR2_X1 i_2196 (.A(n_2477), .B(n_451), .ZN(n_2478));
   INV_X1 i_2197 (.A(n_2478), .ZN(n_2479));
   OR3_X1 i_2198 (.A1(n_2481), .A2(n_2482), .A3(n_2483), .ZN(n_2480));
   NOR2_X1 i_2199 (.A1(n_474), .A2(n_497), .ZN(n_2481));
   NOR2_X1 i_2200 (.A1(n_451), .A2(n_497), .ZN(n_2482));
   NOR2_X1 i_2201 (.A1(n_451), .A2(n_474), .ZN(n_2483));
   XNOR2_X1 i_2202 (.A(n_428), .B(n_405), .ZN(n_2484));
   XNOR2_X1 i_2203 (.A(n_2484), .B(n_382), .ZN(n_2485));
   INV_X1 i_2204 (.A(n_2485), .ZN(n_2486));
   OR3_X1 i_2205 (.A1(n_2488), .A2(n_2489), .A3(n_2490), .ZN(n_2487));
   NOR2_X1 i_2206 (.A1(n_405), .A2(n_428), .ZN(n_2488));
   NOR2_X1 i_2207 (.A1(n_382), .A2(n_428), .ZN(n_2489));
   NOR2_X1 i_2208 (.A1(n_382), .A2(n_405), .ZN(n_2490));
   FA_X1 i_2209 (.A(n_2448), .B(n_2441), .CI(n_2434), .CO(n_2492), .S(n_2491));
   FA_X1 i_2210 (.A(n_2455), .B(n_2486), .CI(n_2479), .CO(n_2494), .S(n_2493));
   FA_X1 i_2211 (.A(n_2472), .B(n_2461), .CI(n_2491), .CO(n_2496), .S(n_2495));
   FA_X1 i_2212 (.A(n_2463), .B(n_2493), .CI(n_2495), .CO(n_2498), .S(n_2497));
   FA_X1 i_2213 (.A(n_2465), .B(n_2467), .CI(n_2497), .CO(n_2500), .S(n_2499));
   XNOR2_X1 i_2214 (.A(n_567), .B(n_544), .ZN(n_2501));
   XNOR2_X1 i_2215 (.A(n_2501), .B(n_521), .ZN(n_2502));
   INV_X1 i_2216 (.A(n_2502), .ZN(n_2503));
   OR3_X1 i_2217 (.A1(n_2505), .A2(n_2506), .A3(n_2507), .ZN(n_2504));
   NOR2_X1 i_2218 (.A1(n_544), .A2(n_567), .ZN(n_2505));
   NOR2_X1 i_2219 (.A1(n_521), .A2(n_567), .ZN(n_2506));
   NOR2_X1 i_2220 (.A1(n_521), .A2(n_544), .ZN(n_2507));
   XNOR2_X1 i_2221 (.A(n_498), .B(n_475), .ZN(n_2508));
   XNOR2_X1 i_2222 (.A(n_2508), .B(n_452), .ZN(n_2509));
   INV_X1 i_2223 (.A(n_2509), .ZN(n_2510));
   OR3_X1 i_2224 (.A1(n_2512), .A2(n_2513), .A3(n_2514), .ZN(n_2511));
   NOR2_X1 i_2225 (.A1(n_475), .A2(n_498), .ZN(n_2512));
   NOR2_X1 i_2226 (.A1(n_452), .A2(n_498), .ZN(n_2513));
   NOR2_X1 i_2227 (.A1(n_452), .A2(n_475), .ZN(n_2514));
   XNOR2_X1 i_2228 (.A(n_429), .B(n_406), .ZN(n_2515));
   XNOR2_X1 i_2229 (.A(n_2515), .B(n_2487), .ZN(n_2516));
   NAND3_X1 i_2230 (.A1(n_2518), .A2(n_2519), .A3(n_2521), .ZN(n_2517));
   OR2_X1 i_2231 (.A1(n_406), .A2(n_429), .ZN(n_2518));
   NAND2_X1 i_2232 (.A1(n_2487), .A2(n_2520), .ZN(n_2519));
   INV_X1 i_2233 (.A(n_429), .ZN(n_2520));
   NAND2_X1 i_2234 (.A1(n_2487), .A2(n_2522), .ZN(n_2521));
   INV_X1 i_2235 (.A(n_406), .ZN(n_2522));
   FA_X1 i_2236 (.A(n_2480), .B(n_2473), .CI(n_2492), .CO(n_2524), .S(n_2523));
   FA_X1 i_2237 (.A(n_2516), .B(n_2510), .CI(n_2503), .CO(n_2526), .S(n_2525));
   FA_X1 i_2238 (.A(n_2523), .B(n_2494), .CI(n_2496), .CO(n_2528), .S(n_2527));
   FA_X1 i_2239 (.A(n_2525), .B(n_2527), .CI(n_2498), .CO(n_2530), .S(n_2529));
   XNOR2_X1 i_2240 (.A(n_568), .B(n_545), .ZN(n_2531));
   XNOR2_X1 i_2241 (.A(n_2531), .B(n_522), .ZN(n_2532));
   INV_X1 i_2242 (.A(n_2532), .ZN(n_2533));
   OR3_X1 i_2243 (.A1(n_2535), .A2(n_2536), .A3(n_2537), .ZN(n_2534));
   NOR2_X1 i_2244 (.A1(n_545), .A2(n_568), .ZN(n_2535));
   NOR2_X1 i_2245 (.A1(n_522), .A2(n_568), .ZN(n_2536));
   NOR2_X1 i_2246 (.A1(n_522), .A2(n_545), .ZN(n_2537));
   XNOR2_X1 i_2247 (.A(n_499), .B(n_476), .ZN(n_2538));
   XNOR2_X1 i_2248 (.A(n_2538), .B(n_453), .ZN(n_2539));
   INV_X1 i_2249 (.A(n_2539), .ZN(n_2540));
   OR3_X1 i_2250 (.A1(n_2542), .A2(n_2543), .A3(n_2544), .ZN(n_2541));
   NOR2_X1 i_2251 (.A1(n_476), .A2(n_499), .ZN(n_2542));
   NOR2_X1 i_2252 (.A1(n_453), .A2(n_499), .ZN(n_2543));
   NOR2_X1 i_2253 (.A1(n_453), .A2(n_476), .ZN(n_2544));
   XNOR2_X1 i_2254 (.A(n_430), .B(n_2511), .ZN(n_2545));
   XNOR2_X1 i_2255 (.A(n_2545), .B(n_2504), .ZN(n_2546));
   INV_X1 i_2256 (.A(n_2546), .ZN(n_2547));
   NAND3_X1 i_2257 (.A1(n_2549), .A2(n_2551), .A3(n_2552), .ZN(n_2548));
   NAND2_X1 i_2258 (.A1(n_2511), .A2(n_2550), .ZN(n_2549));
   INV_X1 i_2259 (.A(n_430), .ZN(n_2550));
   NAND2_X1 i_2260 (.A1(n_2504), .A2(n_2550), .ZN(n_2551));
   NAND2_X1 i_2261 (.A1(n_2504), .A2(n_2511), .ZN(n_2552));
   FA_X1 i_2262 (.A(n_2517), .B(n_2540), .CI(n_2533), .CO(n_2554), .S(n_2553));
   FA_X1 i_2263 (.A(n_2524), .B(n_2547), .CI(n_2526), .CO(n_2556), .S(n_2555));
   FA_X1 i_2264 (.A(n_2553), .B(n_2528), .CI(n_2555), .CO(n_2558), .S(n_2557));
   XNOR2_X1 i_2265 (.A(n_569), .B(n_546), .ZN(n_2559));
   XNOR2_X1 i_2266 (.A(n_2559), .B(n_523), .ZN(n_2560));
   INV_X1 i_2267 (.A(n_2560), .ZN(n_2561));
   OR3_X1 i_2268 (.A1(n_2563), .A2(n_2564), .A3(n_2565), .ZN(n_2562));
   NOR2_X1 i_2269 (.A1(n_546), .A2(n_569), .ZN(n_2563));
   NOR2_X1 i_2270 (.A1(n_523), .A2(n_569), .ZN(n_2564));
   NOR2_X1 i_2271 (.A1(n_523), .A2(n_546), .ZN(n_2565));
   XNOR2_X1 i_2272 (.A(n_500), .B(n_477), .ZN(n_2566));
   XNOR2_X1 i_2273 (.A(n_2566), .B(n_454), .ZN(n_2567));
   INV_X1 i_2274 (.A(n_2567), .ZN(n_2568));
   OR3_X1 i_2275 (.A1(n_2570), .A2(n_2571), .A3(n_2572), .ZN(n_2569));
   NOR2_X1 i_2276 (.A1(n_477), .A2(n_500), .ZN(n_2570));
   NOR2_X1 i_2277 (.A1(n_454), .A2(n_500), .ZN(n_2571));
   NOR2_X1 i_2278 (.A1(n_454), .A2(n_477), .ZN(n_2572));
   FA_X1 i_2279 (.A(n_2541), .B(n_2534), .CI(n_2548), .CO(n_2574), .S(n_2573));
   FA_X1 i_2280 (.A(n_2568), .B(n_2561), .CI(n_2573), .CO(n_2576), .S(n_2575));
   FA_X1 i_2281 (.A(n_2554), .B(n_2556), .CI(n_2575), .CO(n_2578), .S(n_2577));
   XNOR2_X1 i_2282 (.A(n_570), .B(n_547), .ZN(n_2579));
   XNOR2_X1 i_2283 (.A(n_2579), .B(n_524), .ZN(n_2580));
   INV_X1 i_2284 (.A(n_2580), .ZN(n_2581));
   OR3_X1 i_2285 (.A1(n_2583), .A2(n_2584), .A3(n_2585), .ZN(n_2582));
   NOR2_X1 i_2286 (.A1(n_547), .A2(n_570), .ZN(n_2583));
   NOR2_X1 i_2287 (.A1(n_524), .A2(n_570), .ZN(n_2584));
   NOR2_X1 i_2288 (.A1(n_524), .A2(n_547), .ZN(n_2585));
   XNOR2_X1 i_2289 (.A(n_501), .B(n_478), .ZN(n_2586));
   XNOR2_X1 i_2290 (.A(n_2586), .B(n_2569), .ZN(n_2587));
   NAND3_X1 i_2291 (.A1(n_2589), .A2(n_2590), .A3(n_2592), .ZN(n_2588));
   OR2_X1 i_2292 (.A1(n_478), .A2(n_501), .ZN(n_2589));
   NAND2_X1 i_2293 (.A1(n_2569), .A2(n_2591), .ZN(n_2590));
   INV_X1 i_2294 (.A(n_501), .ZN(n_2591));
   NAND2_X1 i_2295 (.A1(n_2569), .A2(n_2593), .ZN(n_2592));
   INV_X1 i_2296 (.A(n_478), .ZN(n_2593));
   FA_X1 i_2297 (.A(n_2562), .B(n_2587), .CI(n_2581), .CO(n_2595), .S(n_2594));
   FA_X1 i_2298 (.A(n_2574), .B(n_2576), .CI(n_2594), .CO(n_2597), .S(n_2596));
   XNOR2_X1 i_2299 (.A(n_571), .B(n_548), .ZN(n_2598));
   XNOR2_X1 i_2300 (.A(n_2598), .B(n_525), .ZN(n_2599));
   INV_X1 i_2301 (.A(n_2599), .ZN(n_2600));
   OR3_X1 i_2302 (.A1(n_2602), .A2(n_2603), .A3(n_2604), .ZN(n_2601));
   NOR2_X1 i_2303 (.A1(n_548), .A2(n_571), .ZN(n_2602));
   NOR2_X1 i_2304 (.A1(n_525), .A2(n_571), .ZN(n_2603));
   NOR2_X1 i_2305 (.A1(n_525), .A2(n_548), .ZN(n_2604));
   XNOR2_X1 i_2306 (.A(n_502), .B(n_2582), .ZN(n_2605));
   XNOR2_X1 i_2307 (.A(n_2605), .B(n_2588), .ZN(n_2606));
   INV_X1 i_2308 (.A(n_2606), .ZN(n_2607));
   NAND3_X1 i_2309 (.A1(n_2609), .A2(n_2611), .A3(n_2612), .ZN(n_2608));
   NAND2_X1 i_2310 (.A1(n_2582), .A2(n_2610), .ZN(n_2609));
   INV_X1 i_2311 (.A(n_502), .ZN(n_2610));
   NAND2_X1 i_2312 (.A1(n_2588), .A2(n_2610), .ZN(n_2611));
   NAND2_X1 i_2313 (.A1(n_2588), .A2(n_2582), .ZN(n_2612));
   FA_X1 i_2314 (.A(n_2600), .B(n_2607), .CI(n_2595), .CO(n_2614), .S(n_2613));
   XNOR2_X1 i_2315 (.A(n_572), .B(n_549), .ZN(n_2615));
   XNOR2_X1 i_2316 (.A(n_2615), .B(n_526), .ZN(n_2616));
   INV_X1 i_2317 (.A(n_2616), .ZN(n_2617));
   OR3_X1 i_2318 (.A1(n_2619), .A2(n_2620), .A3(n_2621), .ZN(n_2618));
   NOR2_X1 i_2319 (.A1(n_549), .A2(n_572), .ZN(n_2619));
   NOR2_X1 i_2320 (.A1(n_526), .A2(n_572), .ZN(n_2620));
   NOR2_X1 i_2321 (.A1(n_526), .A2(n_549), .ZN(n_2621));
   FA_X1 i_2322 (.A(n_2601), .B(n_2617), .CI(n_2608), .CO(n_2623), .S(n_2622));
   XNOR2_X1 i_2323 (.A(n_573), .B(n_550), .ZN(n_2624));
   XNOR2_X1 i_2324 (.A(n_2624), .B(n_2618), .ZN(n_2625));
   NAND3_X1 i_2325 (.A1(n_2627), .A2(n_2628), .A3(n_2630), .ZN(n_2626));
   OR2_X1 i_2326 (.A1(n_550), .A2(n_573), .ZN(n_2627));
   NAND2_X1 i_2327 (.A1(n_2618), .A2(n_2629), .ZN(n_2628));
   INV_X1 i_2328 (.A(n_573), .ZN(n_2629));
   NAND2_X1 i_2329 (.A1(n_2618), .A2(n_2631), .ZN(n_2630));
   INV_X1 i_2330 (.A(n_550), .ZN(n_2631));
   NOR2_X1 i_2331 (.A1(n_0), .A2(n_23), .ZN(n_2632));
   NAND3_X1 i_2332 (.A1(n_2634), .A2(n_2636), .A3(n_2637), .ZN(n_2633));
   NAND2_X1 i_2333 (.A1(n_576), .A2(n_2635), .ZN(n_2634));
   INV_X1 i_2334 (.A(n_1), .ZN(n_2635));
   NAND2_X1 i_2335 (.A1(n_2632), .A2(n_2635), .ZN(n_2636));
   NAND2_X1 i_2336 (.A1(n_2632), .A2(n_576), .ZN(n_2637));
   FA_X1 i_2337 (.A(n_585), .B(n_580), .CI(n_2633), .CO(n_2639), .S(n_2638));
   FA_X1 i_2338 (.A(n_590), .B(n_603), .CI(n_2639), .CO(n_2641), .S(n_2640));
   FA_X1 i_2339 (.A(n_621), .B(n_619), .CI(n_2641), .CO(n_2643), .S(n_2642));
   FA_X1 i_2340 (.A(n_647), .B(n_645), .CI(n_2643), .CO(n_2645), .S(n_2644));
   FA_X1 i_2341 (.A(n_673), .B(n_675), .CI(n_2645), .CO(n_2647), .S(n_2646));
   FA_X1 i_2342 (.A(n_702), .B(n_704), .CI(n_2647), .CO(n_2649), .S(n_2648));
   FA_X1 i_2343 (.A(n_741), .B(n_739), .CI(n_2649), .CO(n_2651), .S(n_2650));
   FA_X1 i_2344 (.A(n_780), .B(n_778), .CI(n_2651), .CO(n_2653), .S(n_2652));
   FA_X1 i_2345 (.A(n_818), .B(n_820), .CI(n_2653), .CO(n_2655), .S(n_2654));
   FA_X1 i_2346 (.A(n_866), .B(n_868), .CI(n_2655), .CO(n_2657), .S(n_2656));
   FA_X1 i_2347 (.A(n_916), .B(n_918), .CI(n_2657), .CO(n_2659), .S(n_2658));
   FA_X1 i_2348 (.A(n_967), .B(n_969), .CI(n_2659), .CO(n_2661), .S(n_2660));
   FA_X1 i_2349 (.A(n_1026), .B(n_1028), .CI(n_2661), .CO(n_2663), .S(n_2662));
   FA_X1 i_2350 (.A(n_1087), .B(n_1089), .CI(n_2663), .CO(n_2665), .S(n_2664));
   FA_X1 i_2351 (.A(n_1149), .B(n_1151), .CI(n_2665), .CO(n_2667), .S(n_2666));
   FA_X1 i_2352 (.A(n_1152), .B(n_1221), .CI(n_2667), .CO(n_2669), .S(n_2668));
   FA_X1 i_2353 (.A(n_1222), .B(n_1293), .CI(n_2669), .CO(n_2671), .S(n_2670));
   FA_X1 i_2354 (.A(n_1364), .B(n_1366), .CI(n_2671), .CO(n_2673), .S(n_2672));
   FA_X1 i_2355 (.A(n_1367), .B(n_1447), .CI(n_2673), .CO(n_2675), .S(n_2674));
   FA_X1 i_2356 (.A(n_1448), .B(n_1530), .CI(n_2675), .CO(n_2677), .S(n_2676));
   FA_X1 i_2357 (.A(n_1531), .B(n_1614), .CI(n_2677), .CO(n_2678), .S(
      mult_res[23]));
   FA_X1 i_2358 (.A(n_1615), .B(n_1699), .CI(n_2678), .CO(n_2679), .S(
      mult_res[24]));
   FA_X1 i_2359 (.A(n_1700), .B(n_1782), .CI(n_2679), .CO(n_2680), .S(
      mult_res[25]));
   FA_X1 i_2360 (.A(n_1783), .B(n_1857), .CI(n_2680), .CO(n_2681), .S(
      mult_res[26]));
   FA_X1 i_2361 (.A(n_1858), .B(n_1931), .CI(n_2681), .CO(n_2682), .S(
      mult_res[27]));
   FA_X1 i_2362 (.A(n_1932), .B(n_2003), .CI(n_2682), .CO(n_2683), .S(
      mult_res[28]));
   FA_X1 i_2363 (.A(n_2004), .B(n_2067), .CI(n_2683), .CO(n_2684), .S(
      mult_res[29]));
   FA_X1 i_2364 (.A(n_2068), .B(n_2130), .CI(n_2684), .CO(n_2685), .S(
      mult_res[30]));
   FA_X1 i_2365 (.A(n_2131), .B(n_2191), .CI(n_2685), .CO(n_2686), .S(
      mult_res[31]));
   FA_X1 i_2366 (.A(n_2192), .B(n_2244), .CI(n_2686), .CO(n_2687), .S(
      mult_res[32]));
   FA_X1 i_2367 (.A(n_2296), .B(n_2245), .CI(n_2687), .CO(n_2688), .S(
      mult_res[33]));
   FA_X1 i_2368 (.A(n_2297), .B(n_2346), .CI(n_2688), .CO(n_2689), .S(
      mult_res[34]));
   FA_X1 i_2369 (.A(n_2347), .B(n_2388), .CI(n_2689), .CO(n_2690), .S(
      mult_res[35]));
   FA_X1 i_2370 (.A(n_2429), .B(n_2389), .CI(n_2690), .CO(n_2691), .S(
      mult_res[36]));
   FA_X1 i_2371 (.A(n_2430), .B(n_2468), .CI(n_2691), .CO(n_2692), .S(
      mult_res[37]));
   FA_X1 i_2372 (.A(n_2469), .B(n_2499), .CI(n_2692), .CO(n_2693), .S(
      mult_res[38]));
   FA_X1 i_2373 (.A(n_2529), .B(n_2500), .CI(n_2693), .CO(n_2694), .S(
      mult_res[39]));
   FA_X1 i_2374 (.A(n_2530), .B(n_2557), .CI(n_2694), .CO(n_2695), .S(
      mult_res[40]));
   FA_X1 i_2375 (.A(n_2577), .B(n_2558), .CI(n_2695), .CO(n_2696), .S(
      mult_res[41]));
   FA_X1 i_2376 (.A(n_2578), .B(n_2596), .CI(n_2696), .CO(n_2697), .S(
      mult_res[42]));
   FA_X1 i_2377 (.A(n_2613), .B(n_2597), .CI(n_2697), .CO(n_2698), .S(
      mult_res[43]));
   FA_X1 i_2378 (.A(n_2614), .B(n_2622), .CI(n_2698), .CO(n_2699), .S(
      mult_res[44]));
   FA_X1 i_2379 (.A(n_2625), .B(n_2623), .CI(n_2699), .CO(n_2700), .S(
      mult_res[45]));
   XNOR2_X1 i_2380 (.A(n_574), .B(n_2626), .ZN(n_2701));
   XNOR2_X1 i_2381 (.A(n_2701), .B(n_2700), .ZN(n_2702));
   INV_X1 i_2382 (.A(n_2702), .ZN(mult_res[46]));
   NAND3_X1 i_2383 (.A1(n_2703), .A2(n_2705), .A3(n_2706), .ZN(mult_res[47]));
   NAND2_X1 i_2384 (.A1(n_2626), .A2(n_2704), .ZN(n_2703));
   INV_X1 i_2385 (.A(n_574), .ZN(n_2704));
   NAND2_X1 i_2386 (.A1(n_2700), .A2(n_2704), .ZN(n_2705));
   NAND2_X1 i_2387 (.A1(n_2700), .A2(n_2626), .ZN(n_2706));
endmodule

module datapath__0_31(p_0, p_1, shamt);
   input [7:0]p_0;
   output [8:0]p_1;
   input [4:0]shamt;

   XNOR2_X1 i_0 (.A(p_0[0]), .B(shamt[0]), .ZN(n_0));
   INV_X1 i_1 (.A(n_0), .ZN(p_1[0]));
   NAND2_X1 i_2 (.A1(shamt[0]), .A2(n_2), .ZN(n_1));
   INV_X1 i_3 (.A(p_0[0]), .ZN(n_2));
   XNOR2_X1 i_4 (.A(p_0[1]), .B(shamt[1]), .ZN(n_3));
   XNOR2_X1 i_5 (.A(n_3), .B(n_1), .ZN(n_4));
   INV_X1 i_6 (.A(n_4), .ZN(p_1[1]));
   NAND3_X1 i_7 (.A1(n_6), .A2(n_8), .A3(n_9), .ZN(n_5));
   NAND2_X1 i_8 (.A1(p_0[1]), .A2(n_7), .ZN(n_6));
   INV_X1 i_9 (.A(shamt[1]), .ZN(n_7));
   NAND2_X1 i_10 (.A1(n_1), .A2(p_0[1]), .ZN(n_8));
   NAND2_X1 i_11 (.A1(n_1), .A2(n_7), .ZN(n_9));
   XNOR2_X1 i_12 (.A(p_0[2]), .B(shamt[2]), .ZN(n_10));
   XNOR2_X1 i_13 (.A(n_10), .B(n_5), .ZN(n_11));
   INV_X1 i_14 (.A(n_11), .ZN(p_1[2]));
   NAND3_X1 i_15 (.A1(n_13), .A2(n_15), .A3(n_16), .ZN(n_12));
   NAND2_X1 i_16 (.A1(p_0[2]), .A2(n_14), .ZN(n_13));
   INV_X1 i_17 (.A(shamt[2]), .ZN(n_14));
   NAND2_X1 i_18 (.A1(n_5), .A2(p_0[2]), .ZN(n_15));
   NAND2_X1 i_19 (.A1(n_5), .A2(n_14), .ZN(n_16));
   XNOR2_X1 i_20 (.A(p_0[3]), .B(shamt[3]), .ZN(n_17));
   XNOR2_X1 i_21 (.A(n_17), .B(n_12), .ZN(n_18));
   INV_X1 i_22 (.A(n_18), .ZN(p_1[3]));
   NAND3_X1 i_23 (.A1(n_20), .A2(n_22), .A3(n_23), .ZN(n_19));
   NAND2_X1 i_24 (.A1(p_0[3]), .A2(n_21), .ZN(n_20));
   INV_X1 i_25 (.A(shamt[3]), .ZN(n_21));
   NAND2_X1 i_26 (.A1(n_12), .A2(p_0[3]), .ZN(n_22));
   NAND2_X1 i_27 (.A1(n_12), .A2(n_21), .ZN(n_23));
   XNOR2_X1 i_28 (.A(p_0[4]), .B(shamt[4]), .ZN(n_24));
   XNOR2_X1 i_29 (.A(n_24), .B(n_19), .ZN(n_25));
   INV_X1 i_30 (.A(n_25), .ZN(p_1[4]));
   NAND3_X1 i_31 (.A1(n_27), .A2(n_29), .A3(n_30), .ZN(n_26));
   NAND2_X1 i_32 (.A1(p_0[4]), .A2(n_28), .ZN(n_27));
   INV_X1 i_33 (.A(shamt[4]), .ZN(n_28));
   NAND2_X1 i_34 (.A1(n_19), .A2(p_0[4]), .ZN(n_29));
   NAND2_X1 i_35 (.A1(n_19), .A2(n_28), .ZN(n_30));
   XNOR2_X1 i_36 (.A(p_0[5]), .B(n_26), .ZN(p_1[5]));
   OR2_X1 i_37 (.A1(p_0[5]), .A2(n_26), .ZN(n_31));
   XNOR2_X1 i_38 (.A(p_0[6]), .B(n_31), .ZN(p_1[6]));
   OR2_X1 i_39 (.A1(p_0[6]), .A2(n_31), .ZN(n_32));
   XNOR2_X1 i_40 (.A(p_0[7]), .B(n_32), .ZN(p_1[7]));
   OR2_X1 i_41 (.A1(p_0[7]), .A2(n_32), .ZN(n_33));
   INV_X1 i_42 (.A(n_33), .ZN(p_1[8]));
endmodule

module datapath__0_32(Eb, mult_res, p_0, E_sum);
   input [7:0]Eb;
   input mult_res;
   input [7:0]p_0;
   output [8:0]E_sum;

   FA_X1 i_0 (.A(mult_res), .B(p_0[0]), .CI(Eb[0]), .CO(n_0), .S(E_sum[0]));
   FA_X1 i_1 (.A(Eb[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(E_sum[1]));
   FA_X1 i_2 (.A(Eb[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(E_sum[2]));
   FA_X1 i_3 (.A(Eb[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(E_sum[3]));
   FA_X1 i_4 (.A(Eb[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(E_sum[4]));
   FA_X1 i_5 (.A(Eb[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(E_sum[5]));
   FA_X1 i_6 (.A(Eb[6]), .B(p_0[6]), .CI(n_5), .CO(n_6), .S(E_sum[6]));
   FA_X1 i_7 (.A(Eb[7]), .B(p_0[7]), .CI(n_6), .CO(E_sum[8]), .S(E_sum[7]));
endmodule

module datapath__0_33(E_sum, p_0);
   input [8:0]E_sum;
   output [9:0]p_0;

   INV_X1 i_0 (.A(E_sum[0]), .ZN(p_0[0]));
   HA_X1 i_1 (.A(E_sum[1]), .B(E_sum[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(E_sum[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(E_sum[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(E_sum[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(E_sum[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(E_sum[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   XNOR2_X1 i_7 (.A(E_sum[7]), .B(n_5), .ZN(p_0[7]));
   OR2_X1 i_8 (.A1(E_sum[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_9 (.A(E_sum[8]), .B(n_6), .ZN(p_0[8]));
   OR2_X1 i_10 (.A1(E_sum[8]), .A2(n_6), .ZN(n_7));
   INV_X1 i_11 (.A(n_7), .ZN(p_0[9]));
endmodule

module datapath__0_36(p_0, E_sum);
   output [7:0]p_0;
   input [7:0]E_sum;

   INV_X1 i_0 (.A(E_sum[0]), .ZN(n_0));
   XNOR2_X1 i_1 (.A(E_sum[1]), .B(n_0), .ZN(p_0[1]));
   NOR2_X1 i_2 (.A1(E_sum[1]), .A2(E_sum[0]), .ZN(n_1));
   XNOR2_X1 i_3 (.A(E_sum[2]), .B(n_1), .ZN(p_0[2]));
   NOR2_X1 i_4 (.A1(E_sum[2]), .A2(n_3), .ZN(n_2));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   XNOR2_X1 i_6 (.A(E_sum[3]), .B(n_2), .ZN(p_0[3]));
   NOR2_X1 i_7 (.A1(E_sum[3]), .A2(n_5), .ZN(n_4));
   INV_X1 i_8 (.A(n_2), .ZN(n_5));
   XNOR2_X1 i_9 (.A(E_sum[4]), .B(n_4), .ZN(p_0[4]));
   NOR2_X1 i_10 (.A1(E_sum[4]), .A2(n_7), .ZN(n_6));
   INV_X1 i_11 (.A(n_4), .ZN(n_7));
   XNOR2_X1 i_12 (.A(E_sum[5]), .B(n_6), .ZN(p_0[5]));
   NOR2_X1 i_13 (.A1(E_sum[5]), .A2(n_9), .ZN(n_8));
   INV_X1 i_14 (.A(n_6), .ZN(n_9));
   XNOR2_X1 i_15 (.A(E_sum[6]), .B(n_8), .ZN(p_0[6]));
   NOR2_X1 i_16 (.A1(E_sum[6]), .A2(n_11), .ZN(n_10));
   INV_X1 i_17 (.A(n_8), .ZN(n_11));
   XNOR2_X1 i_18 (.A(E_sum[7]), .B(n_10), .ZN(n_12));
   INV_X1 i_19 (.A(n_12), .ZN(p_0[7]));
endmodule

module datapath__0_37(p_0, p_1, p_2);
   input [7:0]p_0;
   input [23:0]p_1;
   output [22:0]p_2;

   MUX2_X1 i_0 (.A(p_1[0]), .B(p_1[16]), .S(p_0[4]), .Z(n_0));
   MUX2_X1 i_1 (.A(p_1[1]), .B(p_1[17]), .S(p_0[4]), .Z(n_1));
   MUX2_X1 i_2 (.A(p_1[2]), .B(p_1[18]), .S(p_0[4]), .Z(n_2));
   MUX2_X1 i_3 (.A(p_1[3]), .B(p_1[19]), .S(p_0[4]), .Z(n_3));
   MUX2_X1 i_4 (.A(p_1[4]), .B(p_1[20]), .S(p_0[4]), .Z(n_4));
   MUX2_X1 i_5 (.A(p_1[5]), .B(p_1[21]), .S(p_0[4]), .Z(n_5));
   MUX2_X1 i_6 (.A(p_1[6]), .B(p_1[22]), .S(p_0[4]), .Z(n_6));
   MUX2_X1 i_7 (.A(p_1[7]), .B(p_1[23]), .S(p_0[4]), .Z(n_7));
   NOR2_X1 i_8 (.A1(n_9), .A2(p_0[4]), .ZN(n_8));
   INV_X1 i_9 (.A(p_1[8]), .ZN(n_9));
   NOR2_X1 i_10 (.A1(n_11), .A2(p_0[4]), .ZN(n_10));
   INV_X1 i_11 (.A(p_1[9]), .ZN(n_11));
   NOR2_X1 i_12 (.A1(n_13), .A2(p_0[4]), .ZN(n_12));
   INV_X1 i_13 (.A(p_1[10]), .ZN(n_13));
   NOR2_X1 i_14 (.A1(n_15), .A2(p_0[4]), .ZN(n_14));
   INV_X1 i_15 (.A(p_1[11]), .ZN(n_15));
   NOR2_X1 i_16 (.A1(n_17), .A2(p_0[4]), .ZN(n_16));
   INV_X1 i_17 (.A(p_1[12]), .ZN(n_17));
   NOR2_X1 i_18 (.A1(n_19), .A2(p_0[4]), .ZN(n_18));
   INV_X1 i_19 (.A(p_1[13]), .ZN(n_19));
   NOR2_X1 i_20 (.A1(n_21), .A2(p_0[4]), .ZN(n_20));
   INV_X1 i_21 (.A(p_1[14]), .ZN(n_21));
   NOR2_X1 i_22 (.A1(n_23), .A2(p_0[4]), .ZN(n_22));
   INV_X1 i_23 (.A(p_1[15]), .ZN(n_23));
   NOR2_X1 i_24 (.A1(n_25), .A2(p_0[4]), .ZN(n_24));
   INV_X1 i_25 (.A(p_1[16]), .ZN(n_25));
   NOR2_X1 i_26 (.A1(n_27), .A2(p_0[4]), .ZN(n_26));
   INV_X1 i_27 (.A(p_1[17]), .ZN(n_27));
   NOR2_X1 i_28 (.A1(n_29), .A2(p_0[4]), .ZN(n_28));
   INV_X1 i_29 (.A(p_1[18]), .ZN(n_29));
   NOR2_X1 i_30 (.A1(n_31), .A2(p_0[4]), .ZN(n_30));
   INV_X1 i_31 (.A(p_1[19]), .ZN(n_31));
   NOR2_X1 i_32 (.A1(n_33), .A2(p_0[4]), .ZN(n_32));
   INV_X1 i_33 (.A(p_1[20]), .ZN(n_33));
   NOR2_X1 i_34 (.A1(n_35), .A2(p_0[4]), .ZN(n_34));
   INV_X1 i_35 (.A(p_1[21]), .ZN(n_35));
   NOR2_X1 i_36 (.A1(n_37), .A2(p_0[4]), .ZN(n_36));
   INV_X1 i_37 (.A(p_1[22]), .ZN(n_37));
   NOR2_X1 i_38 (.A1(n_39), .A2(p_0[4]), .ZN(n_38));
   INV_X1 i_39 (.A(p_1[23]), .ZN(n_39));
   MUX2_X1 i_40 (.A(n_0), .B(n_8), .S(p_0[3]), .Z(n_40));
   MUX2_X1 i_41 (.A(n_1), .B(n_10), .S(p_0[3]), .Z(n_41));
   MUX2_X1 i_42 (.A(n_2), .B(n_12), .S(p_0[3]), .Z(n_42));
   MUX2_X1 i_43 (.A(n_3), .B(n_14), .S(p_0[3]), .Z(n_43));
   MUX2_X1 i_44 (.A(n_4), .B(n_16), .S(p_0[3]), .Z(n_44));
   MUX2_X1 i_45 (.A(n_5), .B(n_18), .S(p_0[3]), .Z(n_45));
   MUX2_X1 i_46 (.A(n_6), .B(n_20), .S(p_0[3]), .Z(n_46));
   MUX2_X1 i_47 (.A(n_7), .B(n_22), .S(p_0[3]), .Z(n_47));
   MUX2_X1 i_48 (.A(n_8), .B(n_24), .S(p_0[3]), .Z(n_48));
   MUX2_X1 i_49 (.A(n_10), .B(n_26), .S(p_0[3]), .Z(n_49));
   MUX2_X1 i_50 (.A(n_12), .B(n_28), .S(p_0[3]), .Z(n_50));
   MUX2_X1 i_51 (.A(n_14), .B(n_30), .S(p_0[3]), .Z(n_51));
   MUX2_X1 i_52 (.A(n_16), .B(n_32), .S(p_0[3]), .Z(n_52));
   MUX2_X1 i_53 (.A(n_18), .B(n_34), .S(p_0[3]), .Z(n_53));
   MUX2_X1 i_54 (.A(n_20), .B(n_36), .S(p_0[3]), .Z(n_54));
   MUX2_X1 i_55 (.A(n_22), .B(n_38), .S(p_0[3]), .Z(n_55));
   NOR2_X1 i_56 (.A1(n_57), .A2(p_0[3]), .ZN(n_56));
   INV_X1 i_57 (.A(n_24), .ZN(n_57));
   NOR2_X1 i_58 (.A1(n_59), .A2(p_0[3]), .ZN(n_58));
   INV_X1 i_59 (.A(n_26), .ZN(n_59));
   NOR2_X1 i_60 (.A1(n_61), .A2(p_0[3]), .ZN(n_60));
   INV_X1 i_61 (.A(n_28), .ZN(n_61));
   NOR2_X1 i_62 (.A1(n_63), .A2(p_0[3]), .ZN(n_62));
   INV_X1 i_63 (.A(n_30), .ZN(n_63));
   NOR2_X1 i_64 (.A1(n_65), .A2(p_0[3]), .ZN(n_64));
   INV_X1 i_65 (.A(n_32), .ZN(n_65));
   NOR2_X1 i_66 (.A1(n_67), .A2(p_0[3]), .ZN(n_66));
   INV_X1 i_67 (.A(n_34), .ZN(n_67));
   NOR2_X1 i_68 (.A1(n_69), .A2(p_0[3]), .ZN(n_68));
   INV_X1 i_69 (.A(n_36), .ZN(n_69));
   NOR2_X1 i_70 (.A1(n_71), .A2(p_0[3]), .ZN(n_70));
   INV_X1 i_71 (.A(n_38), .ZN(n_71));
   MUX2_X1 i_72 (.A(n_40), .B(n_44), .S(p_0[2]), .Z(n_72));
   MUX2_X1 i_73 (.A(n_41), .B(n_45), .S(p_0[2]), .Z(n_73));
   MUX2_X1 i_74 (.A(n_42), .B(n_46), .S(p_0[2]), .Z(n_74));
   MUX2_X1 i_75 (.A(n_43), .B(n_47), .S(p_0[2]), .Z(n_75));
   MUX2_X1 i_76 (.A(n_44), .B(n_48), .S(p_0[2]), .Z(n_76));
   MUX2_X1 i_77 (.A(n_45), .B(n_49), .S(p_0[2]), .Z(n_77));
   MUX2_X1 i_78 (.A(n_46), .B(n_50), .S(p_0[2]), .Z(n_78));
   MUX2_X1 i_79 (.A(n_47), .B(n_51), .S(p_0[2]), .Z(n_79));
   MUX2_X1 i_80 (.A(n_48), .B(n_52), .S(p_0[2]), .Z(n_80));
   MUX2_X1 i_81 (.A(n_49), .B(n_53), .S(p_0[2]), .Z(n_81));
   MUX2_X1 i_82 (.A(n_50), .B(n_54), .S(p_0[2]), .Z(n_82));
   MUX2_X1 i_83 (.A(n_51), .B(n_55), .S(p_0[2]), .Z(n_83));
   MUX2_X1 i_84 (.A(n_52), .B(n_56), .S(p_0[2]), .Z(n_84));
   MUX2_X1 i_85 (.A(n_53), .B(n_58), .S(p_0[2]), .Z(n_85));
   MUX2_X1 i_86 (.A(n_54), .B(n_60), .S(p_0[2]), .Z(n_86));
   MUX2_X1 i_87 (.A(n_55), .B(n_62), .S(p_0[2]), .Z(n_87));
   MUX2_X1 i_88 (.A(n_56), .B(n_64), .S(p_0[2]), .Z(n_88));
   MUX2_X1 i_89 (.A(n_58), .B(n_66), .S(p_0[2]), .Z(n_89));
   MUX2_X1 i_90 (.A(n_60), .B(n_68), .S(p_0[2]), .Z(n_90));
   MUX2_X1 i_91 (.A(n_62), .B(n_70), .S(p_0[2]), .Z(n_91));
   NOR2_X1 i_92 (.A1(n_93), .A2(p_0[2]), .ZN(n_92));
   INV_X1 i_93 (.A(n_64), .ZN(n_93));
   NOR2_X1 i_94 (.A1(n_95), .A2(p_0[2]), .ZN(n_94));
   INV_X1 i_95 (.A(n_66), .ZN(n_95));
   NOR2_X1 i_96 (.A1(n_97), .A2(p_0[2]), .ZN(n_96));
   INV_X1 i_97 (.A(n_68), .ZN(n_97));
   NOR2_X1 i_98 (.A1(n_99), .A2(p_0[2]), .ZN(n_98));
   INV_X1 i_99 (.A(n_70), .ZN(n_99));
   MUX2_X1 i_100 (.A(n_72), .B(n_74), .S(p_0[1]), .Z(n_100));
   MUX2_X1 i_101 (.A(n_73), .B(n_75), .S(p_0[1]), .Z(n_101));
   MUX2_X1 i_102 (.A(n_74), .B(n_76), .S(p_0[1]), .Z(n_102));
   MUX2_X1 i_103 (.A(n_75), .B(n_77), .S(p_0[1]), .Z(n_103));
   MUX2_X1 i_104 (.A(n_76), .B(n_78), .S(p_0[1]), .Z(n_104));
   MUX2_X1 i_105 (.A(n_77), .B(n_79), .S(p_0[1]), .Z(n_105));
   MUX2_X1 i_106 (.A(n_78), .B(n_80), .S(p_0[1]), .Z(n_106));
   MUX2_X1 i_107 (.A(n_79), .B(n_81), .S(p_0[1]), .Z(n_107));
   MUX2_X1 i_108 (.A(n_80), .B(n_82), .S(p_0[1]), .Z(n_108));
   MUX2_X1 i_109 (.A(n_81), .B(n_83), .S(p_0[1]), .Z(n_109));
   MUX2_X1 i_110 (.A(n_82), .B(n_84), .S(p_0[1]), .Z(n_110));
   MUX2_X1 i_111 (.A(n_83), .B(n_85), .S(p_0[1]), .Z(n_111));
   MUX2_X1 i_112 (.A(n_84), .B(n_86), .S(p_0[1]), .Z(n_112));
   MUX2_X1 i_113 (.A(n_85), .B(n_87), .S(p_0[1]), .Z(n_113));
   MUX2_X1 i_114 (.A(n_86), .B(n_88), .S(p_0[1]), .Z(n_114));
   MUX2_X1 i_115 (.A(n_87), .B(n_89), .S(p_0[1]), .Z(n_115));
   MUX2_X1 i_116 (.A(n_88), .B(n_90), .S(p_0[1]), .Z(n_116));
   MUX2_X1 i_117 (.A(n_89), .B(n_91), .S(p_0[1]), .Z(n_117));
   MUX2_X1 i_118 (.A(n_90), .B(n_92), .S(p_0[1]), .Z(n_118));
   MUX2_X1 i_119 (.A(n_91), .B(n_94), .S(p_0[1]), .Z(n_119));
   MUX2_X1 i_120 (.A(n_92), .B(n_96), .S(p_0[1]), .Z(n_120));
   MUX2_X1 i_121 (.A(n_94), .B(n_98), .S(p_0[1]), .Z(n_121));
   NOR2_X1 i_122 (.A1(n_123), .A2(p_0[1]), .ZN(n_122));
   INV_X1 i_123 (.A(n_96), .ZN(n_123));
   NOR2_X1 i_124 (.A1(n_125), .A2(p_0[1]), .ZN(n_124));
   INV_X1 i_125 (.A(n_98), .ZN(n_125));
   MUX2_X1 i_126 (.A(n_100), .B(n_101), .S(p_0[0]), .Z(n_126));
   MUX2_X1 i_127 (.A(n_101), .B(n_102), .S(p_0[0]), .Z(n_127));
   MUX2_X1 i_128 (.A(n_102), .B(n_103), .S(p_0[0]), .Z(n_128));
   MUX2_X1 i_129 (.A(n_103), .B(n_104), .S(p_0[0]), .Z(n_129));
   MUX2_X1 i_130 (.A(n_104), .B(n_105), .S(p_0[0]), .Z(n_130));
   MUX2_X1 i_131 (.A(n_105), .B(n_106), .S(p_0[0]), .Z(n_131));
   MUX2_X1 i_132 (.A(n_106), .B(n_107), .S(p_0[0]), .Z(n_132));
   MUX2_X1 i_133 (.A(n_107), .B(n_108), .S(p_0[0]), .Z(n_133));
   MUX2_X1 i_134 (.A(n_108), .B(n_109), .S(p_0[0]), .Z(n_134));
   MUX2_X1 i_135 (.A(n_109), .B(n_110), .S(p_0[0]), .Z(n_135));
   MUX2_X1 i_136 (.A(n_110), .B(n_111), .S(p_0[0]), .Z(n_136));
   MUX2_X1 i_137 (.A(n_111), .B(n_112), .S(p_0[0]), .Z(n_137));
   MUX2_X1 i_138 (.A(n_112), .B(n_113), .S(p_0[0]), .Z(n_138));
   MUX2_X1 i_139 (.A(n_113), .B(n_114), .S(p_0[0]), .Z(n_139));
   MUX2_X1 i_140 (.A(n_114), .B(n_115), .S(p_0[0]), .Z(n_140));
   MUX2_X1 i_141 (.A(n_115), .B(n_116), .S(p_0[0]), .Z(n_141));
   MUX2_X1 i_142 (.A(n_116), .B(n_117), .S(p_0[0]), .Z(n_142));
   MUX2_X1 i_143 (.A(n_117), .B(n_118), .S(p_0[0]), .Z(n_143));
   MUX2_X1 i_144 (.A(n_118), .B(n_119), .S(p_0[0]), .Z(n_144));
   MUX2_X1 i_145 (.A(n_119), .B(n_120), .S(p_0[0]), .Z(n_145));
   MUX2_X1 i_146 (.A(n_120), .B(n_121), .S(p_0[0]), .Z(n_146));
   MUX2_X1 i_147 (.A(n_121), .B(n_122), .S(p_0[0]), .Z(n_147));
   MUX2_X1 i_148 (.A(n_122), .B(n_124), .S(p_0[0]), .Z(n_148));
   NOR3_X1 i_149 (.A1(p_0[5]), .A2(p_0[6]), .A3(p_0[7]), .ZN(n_149));
   AND2_X1 i_150 (.A1(n_148), .A2(n_149), .ZN(p_2[22]));
   AND2_X1 i_151 (.A1(n_147), .A2(n_149), .ZN(p_2[21]));
   AND2_X1 i_152 (.A1(n_146), .A2(n_149), .ZN(p_2[20]));
   AND2_X1 i_153 (.A1(n_145), .A2(n_149), .ZN(p_2[19]));
   AND2_X1 i_154 (.A1(n_144), .A2(n_149), .ZN(p_2[18]));
   AND2_X1 i_155 (.A1(n_143), .A2(n_149), .ZN(p_2[17]));
   AND2_X1 i_156 (.A1(n_142), .A2(n_149), .ZN(p_2[16]));
   AND2_X1 i_157 (.A1(n_141), .A2(n_149), .ZN(p_2[15]));
   AND2_X1 i_158 (.A1(n_140), .A2(n_149), .ZN(p_2[14]));
   AND2_X1 i_159 (.A1(n_139), .A2(n_149), .ZN(p_2[13]));
   AND2_X1 i_160 (.A1(n_138), .A2(n_149), .ZN(p_2[12]));
   AND2_X1 i_161 (.A1(n_137), .A2(n_149), .ZN(p_2[11]));
   AND2_X1 i_162 (.A1(n_136), .A2(n_149), .ZN(p_2[10]));
   AND2_X1 i_163 (.A1(n_135), .A2(n_149), .ZN(p_2[9]));
   AND2_X1 i_164 (.A1(n_134), .A2(n_149), .ZN(p_2[8]));
   AND2_X1 i_165 (.A1(n_133), .A2(n_149), .ZN(p_2[7]));
   AND2_X1 i_166 (.A1(n_132), .A2(n_149), .ZN(p_2[6]));
   AND2_X1 i_167 (.A1(n_131), .A2(n_149), .ZN(p_2[5]));
   AND2_X1 i_168 (.A1(n_130), .A2(n_149), .ZN(p_2[4]));
   AND2_X1 i_169 (.A1(n_129), .A2(n_149), .ZN(p_2[3]));
   AND2_X1 i_170 (.A1(n_128), .A2(n_149), .ZN(p_2[2]));
   AND2_X1 i_171 (.A1(n_127), .A2(n_149), .ZN(p_2[1]));
   AND2_X1 i_172 (.A1(n_126), .A2(n_149), .ZN(p_2[0]));
endmodule

module floating(i_a, i_b, i_clk, o_res);
   input [31:0]i_a;
   input [31:0]i_b;
   input i_clk;
   output [31:0]o_res;

   wire enable;
   wire [2:0]outB;
   wire [2:0]outA;
   wire [31:0]special_res;
   wire [4:0]shamt;
   wire n_0_0_0;
   wire bSubn;
   wire n_0_0;
   wire n_0_1;
   wire n_0_3_0;
   wire aSubn;
   wire n_0_4_0;
   wire n_0_4_1;
   wire n_0_4_2;
   wire [7:0]Eb;
   wire n_0_4_3;
   wire n_0_4_4;
   wire n_0_4_5;
   wire n_0_4_6;
   wire n_0_4_7;
   wire n_0_4_8;
   wire n_0_5_0;
   wire n_0_5_1;
   wire n_0_2;
   wire n_0_5_2;
   wire n_0_3;
   wire n_0_5_3;
   wire n_0_4;
   wire n_0_5_4;
   wire n_0_5;
   wire n_0_5_5;
   wire n_0_6;
   wire n_0_5_6;
   wire n_0_7;
   wire n_0_5_7;
   wire n_0_8;
   wire n_0_5_8;
   wire n_0_9;
   wire n_0_5_9;
   wire n_0_10;
   wire n_0_5_10;
   wire n_0_11;
   wire n_0_5_11;
   wire n_0_12;
   wire n_0_5_12;
   wire n_0_13;
   wire n_0_5_13;
   wire n_0_14;
   wire n_0_5_14;
   wire n_0_15;
   wire n_0_5_15;
   wire n_0_16;
   wire n_0_5_16;
   wire n_0_17;
   wire n_0_5_17;
   wire n_0_18;
   wire n_0_5_18;
   wire n_0_19;
   wire n_0_5_19;
   wire n_0_20;
   wire n_0_5_20;
   wire n_0_21;
   wire n_0_5_21;
   wire n_0_22;
   wire n_0_5_22;
   wire n_0_23;
   wire n_0_5_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_5_24;
   wire [23:0]Nb;
   wire n_0_7_0;
   wire n_0_7_1;
   wire [23:0]Na;
   wire n_0_7_2;
   wire n_0_7_3;
   wire n_0_7_4;
   wire n_0_7_5;
   wire n_0_7_6;
   wire n_0_7_7;
   wire n_0_7_8;
   wire n_0_7_9;
   wire n_0_7_10;
   wire n_0_7_11;
   wire n_0_7_12;
   wire n_0_7_13;
   wire n_0_7_14;
   wire n_0_7_15;
   wire n_0_7_16;
   wire n_0_7_17;
   wire n_0_7_18;
   wire n_0_7_19;
   wire n_0_7_20;
   wire n_0_7_21;
   wire n_0_7_22;
   wire n_0_7_23;
   wire n_0_7_24;
   wire [47:0]mult_res;
   wire n_0_9_0;
   wire n_0_9_1;
   wire n_0_26;
   wire n_0_9_2;
   wire n_0_27;
   wire n_0_9_3;
   wire n_0_28;
   wire n_0_9_4;
   wire n_0_29;
   wire n_0_9_5;
   wire n_0_30;
   wire n_0_9_6;
   wire n_0_31;
   wire n_0_9_7;
   wire n_0_32;
   wire n_0_9_8;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire zero;
   wire [8:0]E_sum;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_14_0;
   wire n_0_14_1;
   wire n_0_14_2;
   wire n_0_14_3;
   wire n_0_53;
   wire n_0_14_4;
   wire n_0_54;
   wire n_0_14_5;
   wire n_0_55;
   wire n_0_14_6;
   wire n_0_56;
   wire n_0_14_7;
   wire n_0_57;
   wire n_0_14_8;
   wire n_0_58;
   wire n_0_14_9;
   wire n_0_59;
   wire n_0_14_10;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_17_0;
   wire n_0_17_1;
   wire n_0_17_2;
   wire n_0_91;
   wire n_0_18_0;
   wire n_0_18_1;
   wire n_0_18_2;
   wire n_0_18_3;
   wire n_0_18_4;
   wire n_0_92;
   wire n_0_93;
   wire n_0_18_5;
   wire n_0_94;
   wire n_0_19_0;
   wire [31:0]float_res;
   wire n_0_19_1;
   wire n_0_19_2;
   wire n_0_19_3;
   wire n_0_19_4;
   wire n_0_19_5;
   wire n_0_19_6;
   wire n_0_19_7;
   wire n_0_19_8;
   wire n_0_19_9;
   wire n_0_19_10;
   wire n_0_19_11;
   wire n_0_19_12;
   wire n_0_19_13;
   wire n_0_19_14;
   wire n_0_19_15;
   wire n_0_19_16;
   wire n_0_19_17;
   wire n_0_19_18;
   wire n_0_19_19;
   wire n_0_19_20;
   wire n_0_19_21;
   wire n_0_19_22;
   wire n_0_19_23;
   wire n_0_19_24;
   wire n_0_19_25;
   wire n_0_19_26;
   wire n_0_19_27;
   wire n_0_19_28;
   wire n_0_19_29;
   wire n_0_19_30;
   wire n_0_19_31;
   wire n_0_19_32;
   wire n_0_19_33;
   wire n_0_19_34;
   wire n_0_19_35;
   wire n_0_19_36;
   wire n_0_19_37;
   wire n_0_19_38;
   wire n_0_19_39;
   wire n_0_19_40;
   wire n_0_19_41;
   wire n_0_19_42;
   wire n_0_19_43;
   wire n_0_19_44;
   wire n_0_19_45;
   wire n_0_19_46;
   wire n_0_20_0;
   wire n_0_20_1;
   wire [31:0]res;
   wire n_0_20_2;
   wire n_0_20_3;
   wire n_0_20_4;
   wire n_0_20_5;
   wire n_0_20_6;
   wire n_0_20_7;
   wire n_0_20_8;
   wire n_0_20_9;
   wire n_0_20_10;
   wire n_0_20_11;
   wire n_0_20_12;
   wire n_0_20_13;
   wire n_0_20_14;
   wire n_0_20_15;
   wire n_0_20_16;
   wire n_0_20_17;
   wire n_0_20_18;
   wire n_0_20_19;
   wire n_0_20_20;
   wire n_0_20_21;
   wire n_0_20_22;
   wire n_0_20_23;
   wire n_0_20_24;
   wire n_0_20_25;
   wire n_0_20_26;
   wire n_0_20_27;
   wire n_0_20_28;
   wire n_0_20_29;
   wire n_0_20_30;
   wire n_0_20_31;
   wire n_0_20_32;
   wire Sb;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire b;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire Sa;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;

   n_case ncase (.A({Sa, n_0_125, n_0_126, n_0_127, n_0_128, n_0_129, n_0_130, 
      n_0_131, n_0_132, n_0_133, n_0_134, n_0_135, n_0_136, n_0_137, n_0_138, 
      n_0_139, n_0_140, n_0_141, n_0_142, n_0_143, n_0_144, n_0_145, n_0_146, 
      n_0_147, n_0_148, n_0_149, n_0_150, n_0_151, n_0_152, n_0_153, n_0_154, 
      n_0_155}), .B({Sb, n_0_95, n_0_96, n_0_97, n_0_98, n_0_99, n_0_100, 
      n_0_101, b, n_0_102, n_0_103, n_0_104, n_0_105, n_0_106, n_0_107, n_0_108, 
      n_0_109, n_0_110, n_0_111, n_0_112, n_0_113, n_0_114, n_0_115, n_0_116, 
      n_0_117, n_0_118, n_0_119, n_0_120, n_0_121, n_0_122, n_0_123, n_0_124}), 
      .S(special_res), .outA(outA), .outB(outB), .enable(enable));
   zero_counter zcn (.M({n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, 
      n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2}), .Zcount(shamt));
   INV_X1 i_0_0_0 (.A(outB[0]), .ZN(n_0_0_0));
   NOR3_X1 i_0_0_1 (.A1(n_0_0_0), .A2(outB[1]), .A3(outB[2]), .ZN(bSubn));
   INV_X1 i_0_1_0 (.A(bSubn), .ZN(n_0_0));
   OR2_X1 i_0_2_0 (.A1(b), .A2(bSubn), .ZN(n_0_1));
   INV_X1 i_0_3_0 (.A(outA[0]), .ZN(n_0_3_0));
   NOR3_X1 i_0_3_1 (.A1(n_0_3_0), .A2(outA[1]), .A3(outA[2]), .ZN(aSubn));
   INV_X1 i_0_4_0 (.A(aSubn), .ZN(n_0_4_0));
   INV_X1 i_0_4_1 (.A(n_0_1), .ZN(n_0_4_1));
   AOI22_X1 i_0_4_2 (.A1(n_0_4_0), .A2(n_0_101), .B1(aSubn), .B2(n_0_131), 
      .ZN(n_0_4_2));
   INV_X1 i_0_4_3 (.A(n_0_4_2), .ZN(Eb[1]));
   AOI22_X1 i_0_4_4 (.A1(n_0_4_0), .A2(n_0_100), .B1(aSubn), .B2(n_0_130), 
      .ZN(n_0_4_3));
   INV_X1 i_0_4_5 (.A(n_0_4_3), .ZN(Eb[2]));
   AOI22_X1 i_0_4_6 (.A1(n_0_4_0), .A2(n_0_99), .B1(aSubn), .B2(n_0_129), 
      .ZN(n_0_4_4));
   INV_X1 i_0_4_7 (.A(n_0_4_4), .ZN(Eb[3]));
   AOI22_X1 i_0_4_8 (.A1(n_0_4_0), .A2(n_0_98), .B1(aSubn), .B2(n_0_128), 
      .ZN(n_0_4_5));
   INV_X1 i_0_4_9 (.A(n_0_4_5), .ZN(Eb[4]));
   AOI22_X1 i_0_4_10 (.A1(n_0_4_0), .A2(n_0_97), .B1(aSubn), .B2(n_0_127), 
      .ZN(n_0_4_6));
   INV_X1 i_0_4_11 (.A(n_0_4_6), .ZN(Eb[5]));
   AOI22_X1 i_0_4_12 (.A1(n_0_4_0), .A2(n_0_96), .B1(aSubn), .B2(n_0_126), 
      .ZN(n_0_4_7));
   INV_X1 i_0_4_13 (.A(n_0_4_7), .ZN(Eb[6]));
   AOI22_X1 i_0_4_14 (.A1(n_0_4_0), .A2(n_0_95), .B1(aSubn), .B2(n_0_125), 
      .ZN(n_0_4_8));
   INV_X1 i_0_4_15 (.A(n_0_4_8), .ZN(Eb[7]));
   NAND2_X1 i_0_4_16 (.A1(n_0_4_1), .A2(n_0_4_0), .ZN(Eb[0]));
   INV_X1 i_0_5_0 (.A(aSubn), .ZN(n_0_5_0));
   AOI22_X1 i_0_5_1 (.A1(n_0_5_0), .A2(n_0_124), .B1(n_0_155), .B2(aSubn), 
      .ZN(n_0_5_1));
   INV_X1 i_0_5_2 (.A(n_0_5_1), .ZN(n_0_2));
   AOI22_X1 i_0_5_3 (.A1(n_0_5_0), .A2(n_0_123), .B1(aSubn), .B2(n_0_154), 
      .ZN(n_0_5_2));
   INV_X1 i_0_5_4 (.A(n_0_5_2), .ZN(n_0_3));
   AOI22_X1 i_0_5_5 (.A1(n_0_5_0), .A2(n_0_122), .B1(aSubn), .B2(n_0_153), 
      .ZN(n_0_5_3));
   INV_X1 i_0_5_6 (.A(n_0_5_3), .ZN(n_0_4));
   AOI22_X1 i_0_5_7 (.A1(n_0_5_0), .A2(n_0_121), .B1(aSubn), .B2(n_0_152), 
      .ZN(n_0_5_4));
   INV_X1 i_0_5_8 (.A(n_0_5_4), .ZN(n_0_5));
   AOI22_X1 i_0_5_9 (.A1(n_0_5_0), .A2(n_0_120), .B1(aSubn), .B2(n_0_151), 
      .ZN(n_0_5_5));
   INV_X1 i_0_5_10 (.A(n_0_5_5), .ZN(n_0_6));
   AOI22_X1 i_0_5_11 (.A1(n_0_5_0), .A2(n_0_119), .B1(aSubn), .B2(n_0_150), 
      .ZN(n_0_5_6));
   INV_X1 i_0_5_12 (.A(n_0_5_6), .ZN(n_0_7));
   AOI22_X1 i_0_5_13 (.A1(n_0_5_0), .A2(n_0_118), .B1(aSubn), .B2(n_0_149), 
      .ZN(n_0_5_7));
   INV_X1 i_0_5_14 (.A(n_0_5_7), .ZN(n_0_8));
   AOI22_X1 i_0_5_15 (.A1(n_0_5_0), .A2(n_0_117), .B1(aSubn), .B2(n_0_148), 
      .ZN(n_0_5_8));
   INV_X1 i_0_5_16 (.A(n_0_5_8), .ZN(n_0_9));
   AOI22_X1 i_0_5_17 (.A1(n_0_5_0), .A2(n_0_116), .B1(aSubn), .B2(n_0_147), 
      .ZN(n_0_5_9));
   INV_X1 i_0_5_18 (.A(n_0_5_9), .ZN(n_0_10));
   AOI22_X1 i_0_5_19 (.A1(n_0_5_0), .A2(n_0_115), .B1(aSubn), .B2(n_0_146), 
      .ZN(n_0_5_10));
   INV_X1 i_0_5_20 (.A(n_0_5_10), .ZN(n_0_11));
   AOI22_X1 i_0_5_21 (.A1(n_0_5_0), .A2(n_0_114), .B1(aSubn), .B2(n_0_145), 
      .ZN(n_0_5_11));
   INV_X1 i_0_5_22 (.A(n_0_5_11), .ZN(n_0_12));
   AOI22_X1 i_0_5_23 (.A1(n_0_5_0), .A2(n_0_113), .B1(aSubn), .B2(n_0_144), 
      .ZN(n_0_5_12));
   INV_X1 i_0_5_24 (.A(n_0_5_12), .ZN(n_0_13));
   AOI22_X1 i_0_5_25 (.A1(n_0_5_0), .A2(n_0_112), .B1(aSubn), .B2(n_0_143), 
      .ZN(n_0_5_13));
   INV_X1 i_0_5_26 (.A(n_0_5_13), .ZN(n_0_14));
   AOI22_X1 i_0_5_27 (.A1(n_0_5_0), .A2(n_0_111), .B1(aSubn), .B2(n_0_142), 
      .ZN(n_0_5_14));
   INV_X1 i_0_5_28 (.A(n_0_5_14), .ZN(n_0_15));
   AOI22_X1 i_0_5_29 (.A1(n_0_5_0), .A2(n_0_110), .B1(aSubn), .B2(n_0_141), 
      .ZN(n_0_5_15));
   INV_X1 i_0_5_30 (.A(n_0_5_15), .ZN(n_0_16));
   AOI22_X1 i_0_5_31 (.A1(n_0_5_0), .A2(n_0_109), .B1(aSubn), .B2(n_0_140), 
      .ZN(n_0_5_16));
   INV_X1 i_0_5_32 (.A(n_0_5_16), .ZN(n_0_17));
   AOI22_X1 i_0_5_33 (.A1(n_0_5_0), .A2(n_0_108), .B1(aSubn), .B2(n_0_139), 
      .ZN(n_0_5_17));
   INV_X1 i_0_5_34 (.A(n_0_5_17), .ZN(n_0_18));
   AOI22_X1 i_0_5_35 (.A1(n_0_5_0), .A2(n_0_107), .B1(aSubn), .B2(n_0_138), 
      .ZN(n_0_5_18));
   INV_X1 i_0_5_36 (.A(n_0_5_18), .ZN(n_0_19));
   AOI22_X1 i_0_5_37 (.A1(n_0_5_0), .A2(n_0_106), .B1(aSubn), .B2(n_0_137), 
      .ZN(n_0_5_19));
   INV_X1 i_0_5_38 (.A(n_0_5_19), .ZN(n_0_20));
   AOI22_X1 i_0_5_39 (.A1(n_0_5_0), .A2(n_0_105), .B1(aSubn), .B2(n_0_136), 
      .ZN(n_0_5_20));
   INV_X1 i_0_5_40 (.A(n_0_5_20), .ZN(n_0_21));
   AOI22_X1 i_0_5_41 (.A1(n_0_5_0), .A2(n_0_104), .B1(aSubn), .B2(n_0_135), 
      .ZN(n_0_5_21));
   INV_X1 i_0_5_42 (.A(n_0_5_21), .ZN(n_0_22));
   AOI22_X1 i_0_5_43 (.A1(n_0_5_0), .A2(n_0_103), .B1(aSubn), .B2(n_0_134), 
      .ZN(n_0_5_22));
   INV_X1 i_0_5_44 (.A(n_0_5_22), .ZN(n_0_23));
   AOI22_X1 i_0_5_45 (.A1(n_0_5_0), .A2(n_0_102), .B1(aSubn), .B2(n_0_133), 
      .ZN(n_0_5_23));
   INV_X1 i_0_5_46 (.A(n_0_5_23), .ZN(n_0_24));
   INV_X1 i_0_5_47 (.A(n_0_5_24), .ZN(n_0_25));
   NAND2_X1 i_0_5_48 (.A1(n_0_0), .A2(n_0_5_0), .ZN(n_0_5_24));
   datapath i_0_6 (.shamt(shamt), .subn({n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2}), 
      .Nb(Nb));
   INV_X1 i_0_7_0 (.A(aSubn), .ZN(n_0_7_0));
   AOI22_X1 i_0_7_1 (.A1(n_0_7_0), .A2(n_0_155), .B1(n_0_124), .B2(aSubn), 
      .ZN(n_0_7_1));
   INV_X1 i_0_7_2 (.A(n_0_7_1), .ZN(Na[0]));
   AOI22_X1 i_0_7_3 (.A1(n_0_7_0), .A2(n_0_154), .B1(aSubn), .B2(n_0_123), 
      .ZN(n_0_7_2));
   INV_X1 i_0_7_4 (.A(n_0_7_2), .ZN(Na[1]));
   AOI22_X1 i_0_7_5 (.A1(n_0_7_0), .A2(n_0_153), .B1(aSubn), .B2(n_0_122), 
      .ZN(n_0_7_3));
   INV_X1 i_0_7_6 (.A(n_0_7_3), .ZN(Na[2]));
   AOI22_X1 i_0_7_7 (.A1(n_0_7_0), .A2(n_0_152), .B1(aSubn), .B2(n_0_121), 
      .ZN(n_0_7_4));
   INV_X1 i_0_7_8 (.A(n_0_7_4), .ZN(Na[3]));
   AOI22_X1 i_0_7_9 (.A1(n_0_7_0), .A2(n_0_151), .B1(aSubn), .B2(n_0_120), 
      .ZN(n_0_7_5));
   INV_X1 i_0_7_10 (.A(n_0_7_5), .ZN(Na[4]));
   AOI22_X1 i_0_7_11 (.A1(n_0_7_0), .A2(n_0_150), .B1(aSubn), .B2(n_0_119), 
      .ZN(n_0_7_6));
   INV_X1 i_0_7_12 (.A(n_0_7_6), .ZN(Na[5]));
   AOI22_X1 i_0_7_13 (.A1(n_0_7_0), .A2(n_0_149), .B1(aSubn), .B2(n_0_118), 
      .ZN(n_0_7_7));
   INV_X1 i_0_7_14 (.A(n_0_7_7), .ZN(Na[6]));
   AOI22_X1 i_0_7_15 (.A1(n_0_7_0), .A2(n_0_148), .B1(aSubn), .B2(n_0_117), 
      .ZN(n_0_7_8));
   INV_X1 i_0_7_16 (.A(n_0_7_8), .ZN(Na[7]));
   AOI22_X1 i_0_7_17 (.A1(n_0_7_0), .A2(n_0_147), .B1(aSubn), .B2(n_0_116), 
      .ZN(n_0_7_9));
   INV_X1 i_0_7_18 (.A(n_0_7_9), .ZN(Na[8]));
   AOI22_X1 i_0_7_19 (.A1(n_0_7_0), .A2(n_0_146), .B1(aSubn), .B2(n_0_115), 
      .ZN(n_0_7_10));
   INV_X1 i_0_7_20 (.A(n_0_7_10), .ZN(Na[9]));
   AOI22_X1 i_0_7_21 (.A1(n_0_7_0), .A2(n_0_145), .B1(aSubn), .B2(n_0_114), 
      .ZN(n_0_7_11));
   INV_X1 i_0_7_22 (.A(n_0_7_11), .ZN(Na[10]));
   AOI22_X1 i_0_7_23 (.A1(n_0_7_0), .A2(n_0_144), .B1(aSubn), .B2(n_0_113), 
      .ZN(n_0_7_12));
   INV_X1 i_0_7_24 (.A(n_0_7_12), .ZN(Na[11]));
   AOI22_X1 i_0_7_25 (.A1(n_0_7_0), .A2(n_0_143), .B1(aSubn), .B2(n_0_112), 
      .ZN(n_0_7_13));
   INV_X1 i_0_7_26 (.A(n_0_7_13), .ZN(Na[12]));
   AOI22_X1 i_0_7_27 (.A1(n_0_7_0), .A2(n_0_142), .B1(aSubn), .B2(n_0_111), 
      .ZN(n_0_7_14));
   INV_X1 i_0_7_28 (.A(n_0_7_14), .ZN(Na[13]));
   AOI22_X1 i_0_7_29 (.A1(n_0_7_0), .A2(n_0_141), .B1(aSubn), .B2(n_0_110), 
      .ZN(n_0_7_15));
   INV_X1 i_0_7_30 (.A(n_0_7_15), .ZN(Na[14]));
   AOI22_X1 i_0_7_31 (.A1(n_0_7_0), .A2(n_0_140), .B1(aSubn), .B2(n_0_109), 
      .ZN(n_0_7_16));
   INV_X1 i_0_7_32 (.A(n_0_7_16), .ZN(Na[15]));
   AOI22_X1 i_0_7_33 (.A1(n_0_7_0), .A2(n_0_139), .B1(aSubn), .B2(n_0_108), 
      .ZN(n_0_7_17));
   INV_X1 i_0_7_34 (.A(n_0_7_17), .ZN(Na[16]));
   AOI22_X1 i_0_7_35 (.A1(n_0_7_0), .A2(n_0_138), .B1(aSubn), .B2(n_0_107), 
      .ZN(n_0_7_18));
   INV_X1 i_0_7_36 (.A(n_0_7_18), .ZN(Na[17]));
   AOI22_X1 i_0_7_37 (.A1(n_0_7_0), .A2(n_0_137), .B1(aSubn), .B2(n_0_106), 
      .ZN(n_0_7_19));
   INV_X1 i_0_7_38 (.A(n_0_7_19), .ZN(Na[18]));
   AOI22_X1 i_0_7_39 (.A1(n_0_7_0), .A2(n_0_136), .B1(aSubn), .B2(n_0_105), 
      .ZN(n_0_7_20));
   INV_X1 i_0_7_40 (.A(n_0_7_20), .ZN(Na[19]));
   AOI22_X1 i_0_7_41 (.A1(n_0_7_0), .A2(n_0_135), .B1(aSubn), .B2(n_0_104), 
      .ZN(n_0_7_21));
   INV_X1 i_0_7_42 (.A(n_0_7_21), .ZN(Na[20]));
   AOI22_X1 i_0_7_43 (.A1(n_0_7_0), .A2(n_0_134), .B1(aSubn), .B2(n_0_103), 
      .ZN(n_0_7_22));
   INV_X1 i_0_7_44 (.A(n_0_7_22), .ZN(Na[21]));
   AOI22_X1 i_0_7_45 (.A1(n_0_7_0), .A2(n_0_133), .B1(aSubn), .B2(n_0_102), 
      .ZN(n_0_7_23));
   INV_X1 i_0_7_46 (.A(n_0_7_23), .ZN(Na[22]));
   INV_X1 i_0_7_47 (.A(n_0_7_24), .ZN(Na[23]));
   NOR2_X1 i_0_7_48 (.A1(n_0_0), .A2(n_0_7_0), .ZN(n_0_7_24));
   datapath__0_29 i_0_8 (.Nb(Nb), .Na(Na), .mult_res({mult_res[47], mult_res[46], 
      mult_res[45], mult_res[44], mult_res[43], mult_res[42], mult_res[41], 
      mult_res[40], mult_res[39], mult_res[38], mult_res[37], mult_res[36], 
      mult_res[35], mult_res[34], mult_res[33], mult_res[32], mult_res[31], 
      mult_res[30], mult_res[29], mult_res[28], mult_res[27], mult_res[26], 
      mult_res[25], mult_res[24], mult_res[23], uc_0, uc_1, uc_2, uc_3, uc_4, 
      uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22}));
   INV_X1 i_0_9_0 (.A(aSubn), .ZN(n_0_9_0));
   AOI22_X1 i_0_9_1 (.A1(n_0_9_0), .A2(n_0_132), .B1(n_0_1), .B2(aSubn), 
      .ZN(n_0_9_1));
   INV_X1 i_0_9_2 (.A(n_0_9_1), .ZN(n_0_26));
   AOI22_X1 i_0_9_3 (.A1(n_0_9_0), .A2(n_0_131), .B1(aSubn), .B2(n_0_101), 
      .ZN(n_0_9_2));
   INV_X1 i_0_9_4 (.A(n_0_9_2), .ZN(n_0_27));
   AOI22_X1 i_0_9_5 (.A1(n_0_9_0), .A2(n_0_130), .B1(aSubn), .B2(n_0_100), 
      .ZN(n_0_9_3));
   INV_X1 i_0_9_6 (.A(n_0_9_3), .ZN(n_0_28));
   AOI22_X1 i_0_9_7 (.A1(n_0_9_0), .A2(n_0_129), .B1(aSubn), .B2(n_0_99), 
      .ZN(n_0_9_4));
   INV_X1 i_0_9_8 (.A(n_0_9_4), .ZN(n_0_29));
   AOI22_X1 i_0_9_9 (.A1(n_0_9_0), .A2(n_0_128), .B1(aSubn), .B2(n_0_98), 
      .ZN(n_0_9_5));
   INV_X1 i_0_9_10 (.A(n_0_9_5), .ZN(n_0_30));
   AOI22_X1 i_0_9_11 (.A1(n_0_9_0), .A2(n_0_127), .B1(aSubn), .B2(n_0_97), 
      .ZN(n_0_9_6));
   INV_X1 i_0_9_12 (.A(n_0_9_6), .ZN(n_0_31));
   AOI22_X1 i_0_9_13 (.A1(n_0_9_0), .A2(n_0_126), .B1(aSubn), .B2(n_0_96), 
      .ZN(n_0_9_7));
   INV_X1 i_0_9_14 (.A(n_0_9_7), .ZN(n_0_32));
   AOI22_X1 i_0_9_15 (.A1(n_0_9_0), .A2(n_0_125), .B1(aSubn), .B2(n_0_95), 
      .ZN(n_0_9_8));
   INV_X1 i_0_9_16 (.A(n_0_9_8), .ZN(n_0_33));
   datapath__0_31 i_0_10 (.p_0({n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26}), .p_1({zero, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
      n_0_36, n_0_35, n_0_34}), .shamt(shamt));
   datapath__0_32 i_0_11 (.Eb(Eb), .mult_res(mult_res[47]), .p_0({n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34}), .E_sum(E_sum));
   datapath__0_33 i_0_12 (.E_sum(E_sum), .p_0({n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42}));
   OR2_X1 i_0_13_0 (.A1(n_0_51), .A2(zero), .ZN(n_0_52));
   INV_X1 i_0_14_0 (.A(n_0_52), .ZN(n_0_14_0));
   NAND2_X1 i_0_14_1 (.A1(n_0_14_0), .A2(n_0_50), .ZN(n_0_14_1));
   OR2_X1 i_0_14_2 (.A1(n_0_50), .A2(n_0_52), .ZN(n_0_14_2));
   INV_X1 i_0_14_3 (.A(n_0_42), .ZN(n_0_14_3));
   OAI21_X1 i_0_14_4 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_3), .ZN(n_0_53));
   INV_X1 i_0_14_5 (.A(n_0_43), .ZN(n_0_14_4));
   OAI21_X1 i_0_14_6 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_4), .ZN(n_0_54));
   INV_X1 i_0_14_7 (.A(n_0_44), .ZN(n_0_14_5));
   OAI21_X1 i_0_14_8 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_5), .ZN(n_0_55));
   INV_X1 i_0_14_9 (.A(n_0_45), .ZN(n_0_14_6));
   OAI21_X1 i_0_14_10 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_6), .ZN(n_0_56));
   INV_X1 i_0_14_11 (.A(n_0_46), .ZN(n_0_14_7));
   OAI21_X1 i_0_14_12 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_7), .ZN(n_0_57));
   INV_X1 i_0_14_13 (.A(n_0_47), .ZN(n_0_14_8));
   OAI21_X1 i_0_14_14 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_8), .ZN(n_0_58));
   INV_X1 i_0_14_15 (.A(n_0_48), .ZN(n_0_14_9));
   OAI21_X1 i_0_14_16 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_9), .ZN(n_0_59));
   INV_X1 i_0_14_17 (.A(n_0_49), .ZN(n_0_14_10));
   OAI21_X1 i_0_14_18 (.A(n_0_14_1), .B1(n_0_14_2), .B2(n_0_14_10), .ZN(n_0_60));
   datapath__0_36 i_0_15 (.p_0({n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, 
      n_0_61, uc_23}), .E_sum({E_sum[7], E_sum[6], E_sum[5], E_sum[4], E_sum[3], 
      E_sum[2], E_sum[1], E_sum[0]}));
   datapath__0_37 i_0_16 (.p_0({n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, 
      n_0_61, E_sum[0]}), .p_1({mult_res[46], mult_res[45], mult_res[44], 
      mult_res[43], mult_res[42], mult_res[41], mult_res[40], mult_res[39], 
      mult_res[38], mult_res[37], mult_res[36], mult_res[35], mult_res[34], 
      mult_res[33], mult_res[32], mult_res[31], mult_res[30], mult_res[29], 
      mult_res[28], mult_res[27], mult_res[26], mult_res[25], mult_res[24], 
      mult_res[23]}), .p_2({n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, 
      n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68}));
   AND4_X1 i_0_17_0 (.A1(n_0_57), .A2(n_0_58), .A3(n_0_59), .A4(n_0_60), 
      .ZN(n_0_17_0));
   AND4_X1 i_0_17_1 (.A1(n_0_17_0), .A2(n_0_54), .A3(n_0_55), .A4(n_0_56), 
      .ZN(n_0_17_1));
   AOI21_X1 i_0_17_2 (.A(zero), .B1(n_0_17_1), .B2(n_0_53), .ZN(n_0_17_2));
   INV_X1 i_0_17_3 (.A(n_0_17_2), .ZN(n_0_91));
   NOR4_X1 i_0_18_0 (.A1(n_0_53), .A2(n_0_54), .A3(n_0_55), .A4(n_0_56), 
      .ZN(n_0_18_0));
   NOR4_X1 i_0_18_1 (.A1(n_0_57), .A2(n_0_58), .A3(n_0_59), .A4(n_0_60), 
      .ZN(n_0_18_1));
   NAND2_X1 i_0_18_2 (.A1(n_0_18_0), .A2(n_0_18_1), .ZN(n_0_18_2));
   INV_X1 i_0_18_3 (.A(n_0_91), .ZN(n_0_18_3));
   NAND2_X1 i_0_18_4 (.A1(n_0_18_2), .A2(n_0_18_3), .ZN(n_0_18_4));
   NOR2_X1 i_0_18_5 (.A1(n_0_18_4), .A2(mult_res[47]), .ZN(n_0_92));
   NOR2_X1 i_0_18_6 (.A1(n_0_18_2), .A2(n_0_91), .ZN(n_0_93));
   INV_X1 i_0_18_7 (.A(mult_res[47]), .ZN(n_0_18_5));
   NOR2_X1 i_0_18_8 (.A1(n_0_18_4), .A2(n_0_18_5), .ZN(n_0_94));
   AOI222_X1 i_0_19_0 (.A1(n_0_68), .A2(n_0_93), .B1(mult_res[24]), .B2(n_0_94), 
      .C1(mult_res[23]), .C2(n_0_92), .ZN(n_0_19_0));
   INV_X1 i_0_19_1 (.A(n_0_19_0), .ZN(float_res[0]));
   NAND2_X1 i_0_19_2 (.A1(n_0_93), .A2(n_0_69), .ZN(n_0_19_1));
   INV_X1 i_0_19_3 (.A(n_0_94), .ZN(n_0_19_2));
   INV_X1 i_0_19_4 (.A(mult_res[25]), .ZN(n_0_19_3));
   INV_X1 i_0_19_5 (.A(mult_res[24]), .ZN(n_0_19_4));
   INV_X1 i_0_19_6 (.A(n_0_92), .ZN(n_0_19_5));
   OAI221_X1 i_0_19_7 (.A(n_0_19_1), .B1(n_0_19_2), .B2(n_0_19_3), .C1(n_0_19_4), 
      .C2(n_0_19_5), .ZN(float_res[1]));
   NAND2_X1 i_0_19_8 (.A1(n_0_93), .A2(n_0_70), .ZN(n_0_19_6));
   INV_X1 i_0_19_9 (.A(mult_res[26]), .ZN(n_0_19_7));
   OAI221_X1 i_0_19_10 (.A(n_0_19_6), .B1(n_0_19_2), .B2(n_0_19_7), .C1(n_0_19_5), 
      .C2(n_0_19_3), .ZN(float_res[2]));
   NAND2_X1 i_0_19_11 (.A1(n_0_93), .A2(n_0_71), .ZN(n_0_19_8));
   INV_X1 i_0_19_12 (.A(mult_res[27]), .ZN(n_0_19_9));
   OAI221_X1 i_0_19_13 (.A(n_0_19_8), .B1(n_0_19_2), .B2(n_0_19_9), .C1(n_0_19_5), 
      .C2(n_0_19_7), .ZN(float_res[3]));
   NAND2_X1 i_0_19_14 (.A1(n_0_93), .A2(n_0_72), .ZN(n_0_19_10));
   INV_X1 i_0_19_15 (.A(mult_res[28]), .ZN(n_0_19_11));
   OAI221_X1 i_0_19_16 (.A(n_0_19_10), .B1(n_0_19_2), .B2(n_0_19_11), .C1(
      n_0_19_5), .C2(n_0_19_9), .ZN(float_res[4]));
   NAND2_X1 i_0_19_17 (.A1(n_0_93), .A2(n_0_73), .ZN(n_0_19_12));
   INV_X1 i_0_19_18 (.A(mult_res[29]), .ZN(n_0_19_13));
   OAI221_X1 i_0_19_19 (.A(n_0_19_12), .B1(n_0_19_2), .B2(n_0_19_13), .C1(
      n_0_19_5), .C2(n_0_19_11), .ZN(float_res[5]));
   NAND2_X1 i_0_19_20 (.A1(n_0_93), .A2(n_0_74), .ZN(n_0_19_14));
   INV_X1 i_0_19_21 (.A(mult_res[30]), .ZN(n_0_19_15));
   OAI221_X1 i_0_19_22 (.A(n_0_19_14), .B1(n_0_19_2), .B2(n_0_19_15), .C1(
      n_0_19_5), .C2(n_0_19_13), .ZN(float_res[6]));
   NAND2_X1 i_0_19_23 (.A1(n_0_93), .A2(n_0_75), .ZN(n_0_19_16));
   INV_X1 i_0_19_24 (.A(mult_res[31]), .ZN(n_0_19_17));
   OAI221_X1 i_0_19_25 (.A(n_0_19_16), .B1(n_0_19_2), .B2(n_0_19_17), .C1(
      n_0_19_5), .C2(n_0_19_15), .ZN(float_res[7]));
   NAND2_X1 i_0_19_26 (.A1(n_0_93), .A2(n_0_76), .ZN(n_0_19_18));
   INV_X1 i_0_19_27 (.A(mult_res[32]), .ZN(n_0_19_19));
   OAI221_X1 i_0_19_28 (.A(n_0_19_18), .B1(n_0_19_2), .B2(n_0_19_19), .C1(
      n_0_19_5), .C2(n_0_19_17), .ZN(float_res[8]));
   NAND2_X1 i_0_19_29 (.A1(n_0_93), .A2(n_0_77), .ZN(n_0_19_20));
   INV_X1 i_0_19_30 (.A(mult_res[33]), .ZN(n_0_19_21));
   OAI221_X1 i_0_19_31 (.A(n_0_19_20), .B1(n_0_19_2), .B2(n_0_19_21), .C1(
      n_0_19_5), .C2(n_0_19_19), .ZN(float_res[9]));
   NAND2_X1 i_0_19_32 (.A1(n_0_93), .A2(n_0_78), .ZN(n_0_19_22));
   INV_X1 i_0_19_33 (.A(mult_res[34]), .ZN(n_0_19_23));
   OAI221_X1 i_0_19_34 (.A(n_0_19_22), .B1(n_0_19_2), .B2(n_0_19_23), .C1(
      n_0_19_5), .C2(n_0_19_21), .ZN(float_res[10]));
   NAND2_X1 i_0_19_35 (.A1(n_0_93), .A2(n_0_79), .ZN(n_0_19_24));
   INV_X1 i_0_19_36 (.A(mult_res[35]), .ZN(n_0_19_25));
   OAI221_X1 i_0_19_37 (.A(n_0_19_24), .B1(n_0_19_2), .B2(n_0_19_25), .C1(
      n_0_19_5), .C2(n_0_19_23), .ZN(float_res[11]));
   NAND2_X1 i_0_19_38 (.A1(n_0_93), .A2(n_0_80), .ZN(n_0_19_26));
   INV_X1 i_0_19_39 (.A(mult_res[36]), .ZN(n_0_19_27));
   OAI221_X1 i_0_19_40 (.A(n_0_19_26), .B1(n_0_19_2), .B2(n_0_19_27), .C1(
      n_0_19_5), .C2(n_0_19_25), .ZN(float_res[12]));
   NAND2_X1 i_0_19_41 (.A1(n_0_93), .A2(n_0_81), .ZN(n_0_19_28));
   INV_X1 i_0_19_42 (.A(mult_res[37]), .ZN(n_0_19_29));
   OAI221_X1 i_0_19_43 (.A(n_0_19_28), .B1(n_0_19_2), .B2(n_0_19_29), .C1(
      n_0_19_5), .C2(n_0_19_27), .ZN(float_res[13]));
   NAND2_X1 i_0_19_44 (.A1(n_0_93), .A2(n_0_82), .ZN(n_0_19_30));
   INV_X1 i_0_19_45 (.A(mult_res[38]), .ZN(n_0_19_31));
   OAI221_X1 i_0_19_46 (.A(n_0_19_30), .B1(n_0_19_2), .B2(n_0_19_31), .C1(
      n_0_19_5), .C2(n_0_19_29), .ZN(float_res[14]));
   NAND2_X1 i_0_19_47 (.A1(n_0_93), .A2(n_0_83), .ZN(n_0_19_32));
   INV_X1 i_0_19_48 (.A(mult_res[39]), .ZN(n_0_19_33));
   OAI221_X1 i_0_19_49 (.A(n_0_19_32), .B1(n_0_19_2), .B2(n_0_19_33), .C1(
      n_0_19_5), .C2(n_0_19_31), .ZN(float_res[15]));
   NAND2_X1 i_0_19_50 (.A1(n_0_93), .A2(n_0_84), .ZN(n_0_19_34));
   INV_X1 i_0_19_51 (.A(mult_res[40]), .ZN(n_0_19_35));
   OAI221_X1 i_0_19_52 (.A(n_0_19_34), .B1(n_0_19_2), .B2(n_0_19_35), .C1(
      n_0_19_5), .C2(n_0_19_33), .ZN(float_res[16]));
   NAND2_X1 i_0_19_53 (.A1(n_0_93), .A2(n_0_85), .ZN(n_0_19_36));
   INV_X1 i_0_19_54 (.A(mult_res[41]), .ZN(n_0_19_37));
   OAI221_X1 i_0_19_55 (.A(n_0_19_36), .B1(n_0_19_2), .B2(n_0_19_37), .C1(
      n_0_19_5), .C2(n_0_19_35), .ZN(float_res[17]));
   NAND2_X1 i_0_19_56 (.A1(n_0_93), .A2(n_0_86), .ZN(n_0_19_38));
   INV_X1 i_0_19_57 (.A(mult_res[42]), .ZN(n_0_19_39));
   OAI221_X1 i_0_19_58 (.A(n_0_19_38), .B1(n_0_19_2), .B2(n_0_19_39), .C1(
      n_0_19_5), .C2(n_0_19_37), .ZN(float_res[18]));
   NAND2_X1 i_0_19_59 (.A1(n_0_93), .A2(n_0_87), .ZN(n_0_19_40));
   INV_X1 i_0_19_60 (.A(mult_res[43]), .ZN(n_0_19_41));
   OAI221_X1 i_0_19_61 (.A(n_0_19_40), .B1(n_0_19_2), .B2(n_0_19_41), .C1(
      n_0_19_5), .C2(n_0_19_39), .ZN(float_res[19]));
   NAND2_X1 i_0_19_62 (.A1(n_0_93), .A2(n_0_88), .ZN(n_0_19_42));
   INV_X1 i_0_19_63 (.A(mult_res[44]), .ZN(n_0_19_43));
   OAI221_X1 i_0_19_64 (.A(n_0_19_42), .B1(n_0_19_2), .B2(n_0_19_43), .C1(
      n_0_19_5), .C2(n_0_19_41), .ZN(float_res[20]));
   NAND2_X1 i_0_19_65 (.A1(n_0_93), .A2(n_0_89), .ZN(n_0_19_44));
   INV_X1 i_0_19_66 (.A(mult_res[45]), .ZN(n_0_19_45));
   OAI221_X1 i_0_19_67 (.A(n_0_19_44), .B1(n_0_19_2), .B2(n_0_19_45), .C1(
      n_0_19_5), .C2(n_0_19_43), .ZN(float_res[21]));
   AOI222_X1 i_0_19_68 (.A1(n_0_93), .A2(n_0_90), .B1(n_0_94), .B2(mult_res[46]), 
      .C1(n_0_92), .C2(mult_res[45]), .ZN(n_0_19_46));
   INV_X1 i_0_19_69 (.A(n_0_19_46), .ZN(float_res[22]));
   XOR2_X1 i_0_19_70 (.A(Sa), .B(Sb), .Z(float_res[31]));
   INV_X1 i_0_20_0 (.A(enable), .ZN(n_0_20_0));
   AOI22_X1 i_0_20_1 (.A1(n_0_20_0), .A2(special_res[0]), .B1(float_res[0]), 
      .B2(enable), .ZN(n_0_20_1));
   INV_X1 i_0_20_2 (.A(n_0_20_1), .ZN(res[0]));
   AOI22_X1 i_0_20_3 (.A1(n_0_20_0), .A2(special_res[1]), .B1(enable), .B2(
      float_res[1]), .ZN(n_0_20_2));
   INV_X1 i_0_20_4 (.A(n_0_20_2), .ZN(res[1]));
   AOI22_X1 i_0_20_5 (.A1(n_0_20_0), .A2(special_res[2]), .B1(enable), .B2(
      float_res[2]), .ZN(n_0_20_3));
   INV_X1 i_0_20_6 (.A(n_0_20_3), .ZN(res[2]));
   AOI22_X1 i_0_20_7 (.A1(n_0_20_0), .A2(special_res[3]), .B1(enable), .B2(
      float_res[3]), .ZN(n_0_20_4));
   INV_X1 i_0_20_8 (.A(n_0_20_4), .ZN(res[3]));
   AOI22_X1 i_0_20_9 (.A1(n_0_20_0), .A2(special_res[4]), .B1(enable), .B2(
      float_res[4]), .ZN(n_0_20_5));
   INV_X1 i_0_20_10 (.A(n_0_20_5), .ZN(res[4]));
   AOI22_X1 i_0_20_11 (.A1(n_0_20_0), .A2(special_res[5]), .B1(enable), .B2(
      float_res[5]), .ZN(n_0_20_6));
   INV_X1 i_0_20_12 (.A(n_0_20_6), .ZN(res[5]));
   AOI22_X1 i_0_20_13 (.A1(n_0_20_0), .A2(special_res[6]), .B1(enable), .B2(
      float_res[6]), .ZN(n_0_20_7));
   INV_X1 i_0_20_14 (.A(n_0_20_7), .ZN(res[6]));
   AOI22_X1 i_0_20_15 (.A1(n_0_20_0), .A2(special_res[7]), .B1(enable), .B2(
      float_res[7]), .ZN(n_0_20_8));
   INV_X1 i_0_20_16 (.A(n_0_20_8), .ZN(res[7]));
   AOI22_X1 i_0_20_17 (.A1(n_0_20_0), .A2(special_res[8]), .B1(enable), .B2(
      float_res[8]), .ZN(n_0_20_9));
   INV_X1 i_0_20_18 (.A(n_0_20_9), .ZN(res[8]));
   AOI22_X1 i_0_20_19 (.A1(n_0_20_0), .A2(special_res[9]), .B1(enable), .B2(
      float_res[9]), .ZN(n_0_20_10));
   INV_X1 i_0_20_20 (.A(n_0_20_10), .ZN(res[9]));
   AOI22_X1 i_0_20_21 (.A1(n_0_20_0), .A2(special_res[10]), .B1(enable), 
      .B2(float_res[10]), .ZN(n_0_20_11));
   INV_X1 i_0_20_22 (.A(n_0_20_11), .ZN(res[10]));
   AOI22_X1 i_0_20_23 (.A1(n_0_20_0), .A2(special_res[11]), .B1(enable), 
      .B2(float_res[11]), .ZN(n_0_20_12));
   INV_X1 i_0_20_24 (.A(n_0_20_12), .ZN(res[11]));
   AOI22_X1 i_0_20_25 (.A1(n_0_20_0), .A2(special_res[12]), .B1(enable), 
      .B2(float_res[12]), .ZN(n_0_20_13));
   INV_X1 i_0_20_26 (.A(n_0_20_13), .ZN(res[12]));
   AOI22_X1 i_0_20_27 (.A1(n_0_20_0), .A2(special_res[13]), .B1(enable), 
      .B2(float_res[13]), .ZN(n_0_20_14));
   INV_X1 i_0_20_28 (.A(n_0_20_14), .ZN(res[13]));
   AOI22_X1 i_0_20_29 (.A1(n_0_20_0), .A2(special_res[14]), .B1(enable), 
      .B2(float_res[14]), .ZN(n_0_20_15));
   INV_X1 i_0_20_30 (.A(n_0_20_15), .ZN(res[14]));
   AOI22_X1 i_0_20_31 (.A1(n_0_20_0), .A2(special_res[15]), .B1(enable), 
      .B2(float_res[15]), .ZN(n_0_20_16));
   INV_X1 i_0_20_32 (.A(n_0_20_16), .ZN(res[15]));
   AOI22_X1 i_0_20_33 (.A1(n_0_20_0), .A2(special_res[16]), .B1(enable), 
      .B2(float_res[16]), .ZN(n_0_20_17));
   INV_X1 i_0_20_34 (.A(n_0_20_17), .ZN(res[16]));
   AOI22_X1 i_0_20_35 (.A1(n_0_20_0), .A2(special_res[17]), .B1(enable), 
      .B2(float_res[17]), .ZN(n_0_20_18));
   INV_X1 i_0_20_36 (.A(n_0_20_18), .ZN(res[17]));
   AOI22_X1 i_0_20_37 (.A1(n_0_20_0), .A2(special_res[18]), .B1(enable), 
      .B2(float_res[18]), .ZN(n_0_20_19));
   INV_X1 i_0_20_38 (.A(n_0_20_19), .ZN(res[18]));
   AOI22_X1 i_0_20_39 (.A1(n_0_20_0), .A2(special_res[19]), .B1(enable), 
      .B2(float_res[19]), .ZN(n_0_20_20));
   INV_X1 i_0_20_40 (.A(n_0_20_20), .ZN(res[19]));
   AOI22_X1 i_0_20_41 (.A1(n_0_20_0), .A2(special_res[20]), .B1(enable), 
      .B2(float_res[20]), .ZN(n_0_20_21));
   INV_X1 i_0_20_42 (.A(n_0_20_21), .ZN(res[20]));
   AOI22_X1 i_0_20_43 (.A1(n_0_20_0), .A2(special_res[21]), .B1(enable), 
      .B2(float_res[21]), .ZN(n_0_20_22));
   INV_X1 i_0_20_44 (.A(n_0_20_22), .ZN(res[21]));
   AOI22_X1 i_0_20_45 (.A1(n_0_20_0), .A2(special_res[22]), .B1(enable), 
      .B2(float_res[22]), .ZN(n_0_20_23));
   INV_X1 i_0_20_46 (.A(n_0_20_23), .ZN(res[22]));
   AOI22_X1 i_0_20_47 (.A1(n_0_20_0), .A2(special_res[23]), .B1(enable), 
      .B2(n_0_53), .ZN(n_0_20_24));
   INV_X1 i_0_20_48 (.A(n_0_20_24), .ZN(res[23]));
   AOI22_X1 i_0_20_49 (.A1(n_0_20_0), .A2(special_res[24]), .B1(enable), 
      .B2(n_0_54), .ZN(n_0_20_25));
   INV_X1 i_0_20_50 (.A(n_0_20_25), .ZN(res[24]));
   AOI22_X1 i_0_20_51 (.A1(n_0_20_0), .A2(special_res[25]), .B1(enable), 
      .B2(n_0_55), .ZN(n_0_20_26));
   INV_X1 i_0_20_52 (.A(n_0_20_26), .ZN(res[25]));
   AOI22_X1 i_0_20_53 (.A1(n_0_20_0), .A2(special_res[26]), .B1(enable), 
      .B2(n_0_56), .ZN(n_0_20_27));
   INV_X1 i_0_20_54 (.A(n_0_20_27), .ZN(res[26]));
   AOI22_X1 i_0_20_55 (.A1(n_0_20_0), .A2(special_res[27]), .B1(enable), 
      .B2(n_0_57), .ZN(n_0_20_28));
   INV_X1 i_0_20_56 (.A(n_0_20_28), .ZN(res[27]));
   AOI22_X1 i_0_20_57 (.A1(n_0_20_0), .A2(special_res[28]), .B1(enable), 
      .B2(n_0_58), .ZN(n_0_20_29));
   INV_X1 i_0_20_58 (.A(n_0_20_29), .ZN(res[28]));
   AOI22_X1 i_0_20_59 (.A1(n_0_20_0), .A2(special_res[29]), .B1(enable), 
      .B2(n_0_59), .ZN(n_0_20_30));
   INV_X1 i_0_20_60 (.A(n_0_20_30), .ZN(res[29]));
   AOI22_X1 i_0_20_61 (.A1(n_0_20_0), .A2(special_res[30]), .B1(enable), 
      .B2(n_0_60), .ZN(n_0_20_31));
   INV_X1 i_0_20_62 (.A(n_0_20_31), .ZN(res[30]));
   AOI22_X1 i_0_20_63 (.A1(n_0_20_0), .A2(special_res[31]), .B1(enable), 
      .B2(float_res[31]), .ZN(n_0_20_32));
   INV_X1 i_0_20_64 (.A(n_0_20_32), .ZN(res[31]));
   DFF_X1 \o_res_reg[31]  (.D(res[31]), .CK(i_clk), .Q(o_res[31]), .QN());
   DFF_X1 \o_res_reg[30]  (.D(res[30]), .CK(i_clk), .Q(o_res[30]), .QN());
   DFF_X1 \o_res_reg[29]  (.D(res[29]), .CK(i_clk), .Q(o_res[29]), .QN());
   DFF_X1 \o_res_reg[28]  (.D(res[28]), .CK(i_clk), .Q(o_res[28]), .QN());
   DFF_X1 \o_res_reg[27]  (.D(res[27]), .CK(i_clk), .Q(o_res[27]), .QN());
   DFF_X1 \o_res_reg[26]  (.D(res[26]), .CK(i_clk), .Q(o_res[26]), .QN());
   DFF_X1 \o_res_reg[25]  (.D(res[25]), .CK(i_clk), .Q(o_res[25]), .QN());
   DFF_X1 \o_res_reg[24]  (.D(res[24]), .CK(i_clk), .Q(o_res[24]), .QN());
   DFF_X1 \o_res_reg[23]  (.D(res[23]), .CK(i_clk), .Q(o_res[23]), .QN());
   DFF_X1 \o_res_reg[22]  (.D(res[22]), .CK(i_clk), .Q(o_res[22]), .QN());
   DFF_X1 \o_res_reg[21]  (.D(res[21]), .CK(i_clk), .Q(o_res[21]), .QN());
   DFF_X1 \o_res_reg[20]  (.D(res[20]), .CK(i_clk), .Q(o_res[20]), .QN());
   DFF_X1 \o_res_reg[19]  (.D(res[19]), .CK(i_clk), .Q(o_res[19]), .QN());
   DFF_X1 \o_res_reg[18]  (.D(res[18]), .CK(i_clk), .Q(o_res[18]), .QN());
   DFF_X1 \o_res_reg[17]  (.D(res[17]), .CK(i_clk), .Q(o_res[17]), .QN());
   DFF_X1 \o_res_reg[16]  (.D(res[16]), .CK(i_clk), .Q(o_res[16]), .QN());
   DFF_X1 \o_res_reg[15]  (.D(res[15]), .CK(i_clk), .Q(o_res[15]), .QN());
   DFF_X1 \o_res_reg[14]  (.D(res[14]), .CK(i_clk), .Q(o_res[14]), .QN());
   DFF_X1 \o_res_reg[13]  (.D(res[13]), .CK(i_clk), .Q(o_res[13]), .QN());
   DFF_X1 \o_res_reg[12]  (.D(res[12]), .CK(i_clk), .Q(o_res[12]), .QN());
   DFF_X1 \o_res_reg[11]  (.D(res[11]), .CK(i_clk), .Q(o_res[11]), .QN());
   DFF_X1 \o_res_reg[10]  (.D(res[10]), .CK(i_clk), .Q(o_res[10]), .QN());
   DFF_X1 \o_res_reg[9]  (.D(res[9]), .CK(i_clk), .Q(o_res[9]), .QN());
   DFF_X1 \o_res_reg[8]  (.D(res[8]), .CK(i_clk), .Q(o_res[8]), .QN());
   DFF_X1 \o_res_reg[7]  (.D(res[7]), .CK(i_clk), .Q(o_res[7]), .QN());
   DFF_X1 \o_res_reg[6]  (.D(res[6]), .CK(i_clk), .Q(o_res[6]), .QN());
   DFF_X1 \o_res_reg[5]  (.D(res[5]), .CK(i_clk), .Q(o_res[5]), .QN());
   DFF_X1 \o_res_reg[4]  (.D(res[4]), .CK(i_clk), .Q(o_res[4]), .QN());
   DFF_X1 \o_res_reg[3]  (.D(res[3]), .CK(i_clk), .Q(o_res[3]), .QN());
   DFF_X1 \o_res_reg[2]  (.D(res[2]), .CK(i_clk), .Q(o_res[2]), .QN());
   DFF_X1 \o_res_reg[1]  (.D(res[1]), .CK(i_clk), .Q(o_res[1]), .QN());
   DFF_X1 \o_res_reg[0]  (.D(res[0]), .CK(i_clk), .Q(o_res[0]), .QN());
   DFF_X1 \b_reg[31]  (.D(i_b[31]), .CK(i_clk), .Q(Sb), .QN());
   DFF_X1 \b_reg[30]  (.D(i_b[30]), .CK(i_clk), .Q(n_0_95), .QN());
   DFF_X1 \b_reg[29]  (.D(i_b[29]), .CK(i_clk), .Q(n_0_96), .QN());
   DFF_X1 \b_reg[28]  (.D(i_b[28]), .CK(i_clk), .Q(n_0_97), .QN());
   DFF_X1 \b_reg[27]  (.D(i_b[27]), .CK(i_clk), .Q(n_0_98), .QN());
   DFF_X1 \b_reg[26]  (.D(i_b[26]), .CK(i_clk), .Q(n_0_99), .QN());
   DFF_X1 \b_reg[25]  (.D(i_b[25]), .CK(i_clk), .Q(n_0_100), .QN());
   DFF_X1 \b_reg[24]  (.D(i_b[24]), .CK(i_clk), .Q(n_0_101), .QN());
   DFF_X1 \b_reg[23]  (.D(i_b[23]), .CK(i_clk), .Q(b), .QN());
   DFF_X1 \b_reg[22]  (.D(i_b[22]), .CK(i_clk), .Q(n_0_102), .QN());
   DFF_X1 \b_reg[21]  (.D(i_b[21]), .CK(i_clk), .Q(n_0_103), .QN());
   DFF_X1 \b_reg[20]  (.D(i_b[20]), .CK(i_clk), .Q(n_0_104), .QN());
   DFF_X1 \b_reg[19]  (.D(i_b[19]), .CK(i_clk), .Q(n_0_105), .QN());
   DFF_X1 \b_reg[18]  (.D(i_b[18]), .CK(i_clk), .Q(n_0_106), .QN());
   DFF_X1 \b_reg[17]  (.D(i_b[17]), .CK(i_clk), .Q(n_0_107), .QN());
   DFF_X1 \b_reg[16]  (.D(i_b[16]), .CK(i_clk), .Q(n_0_108), .QN());
   DFF_X1 \b_reg[15]  (.D(i_b[15]), .CK(i_clk), .Q(n_0_109), .QN());
   DFF_X1 \b_reg[14]  (.D(i_b[14]), .CK(i_clk), .Q(n_0_110), .QN());
   DFF_X1 \b_reg[13]  (.D(i_b[13]), .CK(i_clk), .Q(n_0_111), .QN());
   DFF_X1 \b_reg[12]  (.D(i_b[12]), .CK(i_clk), .Q(n_0_112), .QN());
   DFF_X1 \b_reg[11]  (.D(i_b[11]), .CK(i_clk), .Q(n_0_113), .QN());
   DFF_X1 \b_reg[10]  (.D(i_b[10]), .CK(i_clk), .Q(n_0_114), .QN());
   DFF_X1 \b_reg[9]  (.D(i_b[9]), .CK(i_clk), .Q(n_0_115), .QN());
   DFF_X1 \b_reg[8]  (.D(i_b[8]), .CK(i_clk), .Q(n_0_116), .QN());
   DFF_X1 \b_reg[7]  (.D(i_b[7]), .CK(i_clk), .Q(n_0_117), .QN());
   DFF_X1 \b_reg[6]  (.D(i_b[6]), .CK(i_clk), .Q(n_0_118), .QN());
   DFF_X1 \b_reg[5]  (.D(i_b[5]), .CK(i_clk), .Q(n_0_119), .QN());
   DFF_X1 \b_reg[4]  (.D(i_b[4]), .CK(i_clk), .Q(n_0_120), .QN());
   DFF_X1 \b_reg[3]  (.D(i_b[3]), .CK(i_clk), .Q(n_0_121), .QN());
   DFF_X1 \b_reg[2]  (.D(i_b[2]), .CK(i_clk), .Q(n_0_122), .QN());
   DFF_X1 \b_reg[1]  (.D(i_b[1]), .CK(i_clk), .Q(n_0_123), .QN());
   DFF_X1 \b_reg[0]  (.D(i_b[0]), .CK(i_clk), .Q(n_0_124), .QN());
   DFF_X1 \a_reg[31]  (.D(i_a[31]), .CK(i_clk), .Q(Sa), .QN());
   DFF_X1 \a_reg[30]  (.D(i_a[30]), .CK(i_clk), .Q(n_0_125), .QN());
   DFF_X1 \a_reg[29]  (.D(i_a[29]), .CK(i_clk), .Q(n_0_126), .QN());
   DFF_X1 \a_reg[28]  (.D(i_a[28]), .CK(i_clk), .Q(n_0_127), .QN());
   DFF_X1 \a_reg[27]  (.D(i_a[27]), .CK(i_clk), .Q(n_0_128), .QN());
   DFF_X1 \a_reg[26]  (.D(i_a[26]), .CK(i_clk), .Q(n_0_129), .QN());
   DFF_X1 \a_reg[25]  (.D(i_a[25]), .CK(i_clk), .Q(n_0_130), .QN());
   DFF_X1 \a_reg[24]  (.D(i_a[24]), .CK(i_clk), .Q(n_0_131), .QN());
   DFF_X1 \a_reg[23]  (.D(i_a[23]), .CK(i_clk), .Q(n_0_132), .QN());
   DFF_X1 \a_reg[22]  (.D(i_a[22]), .CK(i_clk), .Q(n_0_133), .QN());
   DFF_X1 \a_reg[21]  (.D(i_a[21]), .CK(i_clk), .Q(n_0_134), .QN());
   DFF_X1 \a_reg[20]  (.D(i_a[20]), .CK(i_clk), .Q(n_0_135), .QN());
   DFF_X1 \a_reg[19]  (.D(i_a[19]), .CK(i_clk), .Q(n_0_136), .QN());
   DFF_X1 \a_reg[18]  (.D(i_a[18]), .CK(i_clk), .Q(n_0_137), .QN());
   DFF_X1 \a_reg[17]  (.D(i_a[17]), .CK(i_clk), .Q(n_0_138), .QN());
   DFF_X1 \a_reg[16]  (.D(i_a[16]), .CK(i_clk), .Q(n_0_139), .QN());
   DFF_X1 \a_reg[15]  (.D(i_a[15]), .CK(i_clk), .Q(n_0_140), .QN());
   DFF_X1 \a_reg[14]  (.D(i_a[14]), .CK(i_clk), .Q(n_0_141), .QN());
   DFF_X1 \a_reg[13]  (.D(i_a[13]), .CK(i_clk), .Q(n_0_142), .QN());
   DFF_X1 \a_reg[12]  (.D(i_a[12]), .CK(i_clk), .Q(n_0_143), .QN());
   DFF_X1 \a_reg[11]  (.D(i_a[11]), .CK(i_clk), .Q(n_0_144), .QN());
   DFF_X1 \a_reg[10]  (.D(i_a[10]), .CK(i_clk), .Q(n_0_145), .QN());
   DFF_X1 \a_reg[9]  (.D(i_a[9]), .CK(i_clk), .Q(n_0_146), .QN());
   DFF_X1 \a_reg[8]  (.D(i_a[8]), .CK(i_clk), .Q(n_0_147), .QN());
   DFF_X1 \a_reg[7]  (.D(i_a[7]), .CK(i_clk), .Q(n_0_148), .QN());
   DFF_X1 \a_reg[6]  (.D(i_a[6]), .CK(i_clk), .Q(n_0_149), .QN());
   DFF_X1 \a_reg[5]  (.D(i_a[5]), .CK(i_clk), .Q(n_0_150), .QN());
   DFF_X1 \a_reg[4]  (.D(i_a[4]), .CK(i_clk), .Q(n_0_151), .QN());
   DFF_X1 \a_reg[3]  (.D(i_a[3]), .CK(i_clk), .Q(n_0_152), .QN());
   DFF_X1 \a_reg[2]  (.D(i_a[2]), .CK(i_clk), .Q(n_0_153), .QN());
   DFF_X1 \a_reg[1]  (.D(i_a[1]), .CK(i_clk), .Q(n_0_154), .QN());
   DFF_X1 \a_reg[0]  (.D(i_a[0]), .CK(i_clk), .Q(n_0_155), .QN());
endmodule
